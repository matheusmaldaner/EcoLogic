library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity logic_network is
    port (
        inputs : in std_logic_vector(255 downto 0);
        outputs : out std_logic_vector(9 downto 0)
    );
end logic_network;

architecture Behavioral of logic_network is
    signal layer0_outputs : std_logic_vector(2559 downto 0);

begin

    layer0_outputs(0) <= not(inputs(45)) or (inputs(251));
    layer0_outputs(1) <= '1';
    layer0_outputs(2) <= not((inputs(112)) or (inputs(180)));
    layer0_outputs(3) <= not(inputs(200));
    layer0_outputs(4) <= not((inputs(139)) xor (inputs(104)));
    layer0_outputs(5) <= (inputs(227)) or (inputs(251));
    layer0_outputs(6) <= (inputs(242)) xor (inputs(215));
    layer0_outputs(7) <= (inputs(205)) xor (inputs(33));
    layer0_outputs(8) <= not((inputs(61)) or (inputs(42)));
    layer0_outputs(9) <= not(inputs(91)) or (inputs(35));
    layer0_outputs(10) <= inputs(124);
    layer0_outputs(11) <= (inputs(140)) or (inputs(27));
    layer0_outputs(12) <= not(inputs(17)) or (inputs(252));
    layer0_outputs(13) <= not(inputs(59)) or (inputs(239));
    layer0_outputs(14) <= not((inputs(3)) xor (inputs(188)));
    layer0_outputs(15) <= (inputs(228)) or (inputs(49));
    layer0_outputs(16) <= not(inputs(56)) or (inputs(234));
    layer0_outputs(17) <= inputs(159);
    layer0_outputs(18) <= (inputs(128)) xor (inputs(162));
    layer0_outputs(19) <= not((inputs(242)) xor (inputs(7)));
    layer0_outputs(20) <= inputs(0);
    layer0_outputs(21) <= not(inputs(50)) or (inputs(30));
    layer0_outputs(22) <= not((inputs(9)) xor (inputs(86)));
    layer0_outputs(23) <= (inputs(145)) and (inputs(111));
    layer0_outputs(24) <= inputs(189);
    layer0_outputs(25) <= (inputs(147)) and not (inputs(13));
    layer0_outputs(26) <= (inputs(165)) and not (inputs(98));
    layer0_outputs(27) <= (inputs(90)) or (inputs(175));
    layer0_outputs(28) <= not(inputs(101)) or (inputs(0));
    layer0_outputs(29) <= inputs(137);
    layer0_outputs(30) <= (inputs(195)) or (inputs(191));
    layer0_outputs(31) <= inputs(246);
    layer0_outputs(32) <= not((inputs(204)) or (inputs(42)));
    layer0_outputs(33) <= (inputs(187)) or (inputs(110));
    layer0_outputs(34) <= inputs(215);
    layer0_outputs(35) <= (inputs(48)) and not (inputs(129));
    layer0_outputs(36) <= inputs(132);
    layer0_outputs(37) <= not(inputs(94));
    layer0_outputs(38) <= inputs(90);
    layer0_outputs(39) <= (inputs(178)) or (inputs(140));
    layer0_outputs(40) <= not((inputs(225)) xor (inputs(119)));
    layer0_outputs(41) <= (inputs(14)) and not (inputs(9));
    layer0_outputs(42) <= (inputs(168)) and not (inputs(38));
    layer0_outputs(43) <= not(inputs(174));
    layer0_outputs(44) <= (inputs(231)) xor (inputs(250));
    layer0_outputs(45) <= not((inputs(8)) xor (inputs(93)));
    layer0_outputs(46) <= not((inputs(88)) or (inputs(75)));
    layer0_outputs(47) <= not((inputs(153)) and (inputs(197)));
    layer0_outputs(48) <= (inputs(65)) or (inputs(49));
    layer0_outputs(49) <= (inputs(198)) xor (inputs(34));
    layer0_outputs(50) <= not((inputs(193)) or (inputs(76)));
    layer0_outputs(51) <= not((inputs(240)) xor (inputs(228)));
    layer0_outputs(52) <= not(inputs(100)) or (inputs(20));
    layer0_outputs(53) <= (inputs(117)) or (inputs(1));
    layer0_outputs(54) <= (inputs(140)) or (inputs(81));
    layer0_outputs(55) <= not((inputs(137)) or (inputs(247)));
    layer0_outputs(56) <= (inputs(93)) or (inputs(78));
    layer0_outputs(57) <= not(inputs(166));
    layer0_outputs(58) <= not(inputs(205));
    layer0_outputs(59) <= not((inputs(8)) and (inputs(219)));
    layer0_outputs(60) <= (inputs(71)) or (inputs(29));
    layer0_outputs(61) <= inputs(134);
    layer0_outputs(62) <= (inputs(31)) and (inputs(7));
    layer0_outputs(63) <= inputs(119);
    layer0_outputs(64) <= (inputs(54)) xor (inputs(161));
    layer0_outputs(65) <= not((inputs(211)) or (inputs(148)));
    layer0_outputs(66) <= not((inputs(127)) xor (inputs(51)));
    layer0_outputs(67) <= not(inputs(122)) or (inputs(18));
    layer0_outputs(68) <= not((inputs(17)) xor (inputs(237)));
    layer0_outputs(69) <= not(inputs(78));
    layer0_outputs(70) <= not((inputs(41)) or (inputs(180)));
    layer0_outputs(71) <= inputs(199);
    layer0_outputs(72) <= not((inputs(254)) xor (inputs(68)));
    layer0_outputs(73) <= not(inputs(88));
    layer0_outputs(74) <= (inputs(187)) or (inputs(250));
    layer0_outputs(75) <= not((inputs(75)) or (inputs(33)));
    layer0_outputs(76) <= inputs(190);
    layer0_outputs(77) <= not((inputs(97)) xor (inputs(244)));
    layer0_outputs(78) <= inputs(157);
    layer0_outputs(79) <= not((inputs(22)) xor (inputs(178)));
    layer0_outputs(80) <= (inputs(217)) xor (inputs(1));
    layer0_outputs(81) <= inputs(133);
    layer0_outputs(82) <= inputs(181);
    layer0_outputs(83) <= (inputs(8)) xor (inputs(23));
    layer0_outputs(84) <= (inputs(81)) or (inputs(233));
    layer0_outputs(85) <= not((inputs(79)) or (inputs(188)));
    layer0_outputs(86) <= (inputs(106)) and not (inputs(81));
    layer0_outputs(87) <= not((inputs(229)) xor (inputs(19)));
    layer0_outputs(88) <= inputs(102);
    layer0_outputs(89) <= (inputs(24)) xor (inputs(247));
    layer0_outputs(90) <= (inputs(72)) and not (inputs(38));
    layer0_outputs(91) <= '1';
    layer0_outputs(92) <= not((inputs(47)) or (inputs(62)));
    layer0_outputs(93) <= not((inputs(200)) or (inputs(96)));
    layer0_outputs(94) <= not(inputs(56));
    layer0_outputs(95) <= inputs(92);
    layer0_outputs(96) <= not(inputs(13)) or (inputs(89));
    layer0_outputs(97) <= not(inputs(65)) or (inputs(79));
    layer0_outputs(98) <= '1';
    layer0_outputs(99) <= '1';
    layer0_outputs(100) <= (inputs(132)) and not (inputs(113));
    layer0_outputs(101) <= not((inputs(40)) or (inputs(221)));
    layer0_outputs(102) <= inputs(131);
    layer0_outputs(103) <= (inputs(236)) or (inputs(124));
    layer0_outputs(104) <= not((inputs(200)) xor (inputs(209)));
    layer0_outputs(105) <= not((inputs(197)) or (inputs(161)));
    layer0_outputs(106) <= not(inputs(90)) or (inputs(15));
    layer0_outputs(107) <= inputs(235);
    layer0_outputs(108) <= not(inputs(204));
    layer0_outputs(109) <= not((inputs(207)) or (inputs(151)));
    layer0_outputs(110) <= inputs(175);
    layer0_outputs(111) <= not(inputs(187)) or (inputs(110));
    layer0_outputs(112) <= not(inputs(234));
    layer0_outputs(113) <= (inputs(25)) or (inputs(140));
    layer0_outputs(114) <= not((inputs(59)) or (inputs(208)));
    layer0_outputs(115) <= (inputs(247)) or (inputs(162));
    layer0_outputs(116) <= '0';
    layer0_outputs(117) <= not(inputs(138));
    layer0_outputs(118) <= (inputs(4)) xor (inputs(42));
    layer0_outputs(119) <= (inputs(111)) xor (inputs(147));
    layer0_outputs(120) <= not(inputs(101)) or (inputs(173));
    layer0_outputs(121) <= inputs(6);
    layer0_outputs(122) <= not(inputs(181));
    layer0_outputs(123) <= (inputs(149)) and not (inputs(65));
    layer0_outputs(124) <= not(inputs(210)) or (inputs(17));
    layer0_outputs(125) <= (inputs(7)) xor (inputs(149));
    layer0_outputs(126) <= not(inputs(101)) or (inputs(22));
    layer0_outputs(127) <= (inputs(238)) and (inputs(111));
    layer0_outputs(128) <= (inputs(57)) xor (inputs(224));
    layer0_outputs(129) <= not(inputs(147));
    layer0_outputs(130) <= not(inputs(106));
    layer0_outputs(131) <= not(inputs(74)) or (inputs(9));
    layer0_outputs(132) <= '0';
    layer0_outputs(133) <= (inputs(20)) or (inputs(69));
    layer0_outputs(134) <= not(inputs(166)) or (inputs(79));
    layer0_outputs(135) <= (inputs(118)) and not (inputs(146));
    layer0_outputs(136) <= (inputs(184)) xor (inputs(126));
    layer0_outputs(137) <= not((inputs(24)) or (inputs(39)));
    layer0_outputs(138) <= not(inputs(52));
    layer0_outputs(139) <= not((inputs(246)) or (inputs(214)));
    layer0_outputs(140) <= not(inputs(53));
    layer0_outputs(141) <= (inputs(205)) or (inputs(180));
    layer0_outputs(142) <= not((inputs(210)) or (inputs(145)));
    layer0_outputs(143) <= inputs(131);
    layer0_outputs(144) <= not(inputs(222)) or (inputs(216));
    layer0_outputs(145) <= not((inputs(227)) or (inputs(54)));
    layer0_outputs(146) <= (inputs(107)) and not (inputs(13));
    layer0_outputs(147) <= (inputs(255)) and not (inputs(218));
    layer0_outputs(148) <= inputs(138);
    layer0_outputs(149) <= inputs(105);
    layer0_outputs(150) <= (inputs(229)) and not (inputs(47));
    layer0_outputs(151) <= (inputs(94)) xor (inputs(221));
    layer0_outputs(152) <= not(inputs(116));
    layer0_outputs(153) <= not((inputs(193)) xor (inputs(162)));
    layer0_outputs(154) <= not(inputs(211)) or (inputs(46));
    layer0_outputs(155) <= not((inputs(112)) or (inputs(70)));
    layer0_outputs(156) <= not((inputs(138)) and (inputs(17)));
    layer0_outputs(157) <= not(inputs(118));
    layer0_outputs(158) <= not((inputs(136)) or (inputs(11)));
    layer0_outputs(159) <= inputs(166);
    layer0_outputs(160) <= (inputs(187)) or (inputs(45));
    layer0_outputs(161) <= (inputs(69)) or (inputs(187));
    layer0_outputs(162) <= not(inputs(58));
    layer0_outputs(163) <= not((inputs(187)) or (inputs(160)));
    layer0_outputs(164) <= (inputs(155)) and not (inputs(207));
    layer0_outputs(165) <= not(inputs(198));
    layer0_outputs(166) <= inputs(150);
    layer0_outputs(167) <= not((inputs(188)) or (inputs(141)));
    layer0_outputs(168) <= not(inputs(164));
    layer0_outputs(169) <= not((inputs(132)) xor (inputs(82)));
    layer0_outputs(170) <= not(inputs(60));
    layer0_outputs(171) <= (inputs(241)) xor (inputs(21));
    layer0_outputs(172) <= not((inputs(94)) or (inputs(230)));
    layer0_outputs(173) <= (inputs(105)) and not (inputs(237));
    layer0_outputs(174) <= not((inputs(89)) or (inputs(229)));
    layer0_outputs(175) <= not((inputs(208)) or (inputs(183)));
    layer0_outputs(176) <= (inputs(200)) and not (inputs(130));
    layer0_outputs(177) <= (inputs(233)) or (inputs(18));
    layer0_outputs(178) <= not((inputs(59)) or (inputs(230)));
    layer0_outputs(179) <= (inputs(144)) xor (inputs(108));
    layer0_outputs(180) <= (inputs(133)) or (inputs(70));
    layer0_outputs(181) <= not(inputs(81));
    layer0_outputs(182) <= (inputs(6)) or (inputs(148));
    layer0_outputs(183) <= not((inputs(117)) or (inputs(131)));
    layer0_outputs(184) <= not(inputs(104));
    layer0_outputs(185) <= not(inputs(171));
    layer0_outputs(186) <= '0';
    layer0_outputs(187) <= (inputs(174)) or (inputs(181));
    layer0_outputs(188) <= inputs(55);
    layer0_outputs(189) <= not((inputs(159)) and (inputs(9)));
    layer0_outputs(190) <= not((inputs(36)) or (inputs(189)));
    layer0_outputs(191) <= not(inputs(1)) or (inputs(92));
    layer0_outputs(192) <= inputs(231);
    layer0_outputs(193) <= not(inputs(222)) or (inputs(21));
    layer0_outputs(194) <= not((inputs(74)) or (inputs(162)));
    layer0_outputs(195) <= (inputs(199)) and not (inputs(83));
    layer0_outputs(196) <= (inputs(155)) or (inputs(174));
    layer0_outputs(197) <= (inputs(202)) and not (inputs(249));
    layer0_outputs(198) <= (inputs(118)) and not (inputs(229));
    layer0_outputs(199) <= (inputs(110)) and (inputs(66));
    layer0_outputs(200) <= '0';
    layer0_outputs(201) <= not((inputs(84)) or (inputs(163)));
    layer0_outputs(202) <= not(inputs(195)) or (inputs(235));
    layer0_outputs(203) <= inputs(183);
    layer0_outputs(204) <= not((inputs(39)) or (inputs(224)));
    layer0_outputs(205) <= not((inputs(227)) and (inputs(98)));
    layer0_outputs(206) <= inputs(107);
    layer0_outputs(207) <= (inputs(196)) or (inputs(33));
    layer0_outputs(208) <= not((inputs(137)) or (inputs(245)));
    layer0_outputs(209) <= not((inputs(150)) or (inputs(69)));
    layer0_outputs(210) <= inputs(91);
    layer0_outputs(211) <= not((inputs(150)) or (inputs(64)));
    layer0_outputs(212) <= not(inputs(92));
    layer0_outputs(213) <= not(inputs(175)) or (inputs(251));
    layer0_outputs(214) <= not(inputs(152)) or (inputs(154));
    layer0_outputs(215) <= not((inputs(206)) or (inputs(220)));
    layer0_outputs(216) <= inputs(120);
    layer0_outputs(217) <= (inputs(136)) xor (inputs(208));
    layer0_outputs(218) <= not(inputs(90)) or (inputs(56));
    layer0_outputs(219) <= not(inputs(172)) or (inputs(45));
    layer0_outputs(220) <= not((inputs(6)) xor (inputs(139)));
    layer0_outputs(221) <= not(inputs(88)) or (inputs(19));
    layer0_outputs(222) <= not(inputs(245));
    layer0_outputs(223) <= not(inputs(147));
    layer0_outputs(224) <= not((inputs(221)) or (inputs(187)));
    layer0_outputs(225) <= (inputs(195)) or (inputs(69));
    layer0_outputs(226) <= inputs(217);
    layer0_outputs(227) <= not(inputs(133));
    layer0_outputs(228) <= '0';
    layer0_outputs(229) <= inputs(210);
    layer0_outputs(230) <= '0';
    layer0_outputs(231) <= not((inputs(254)) and (inputs(18)));
    layer0_outputs(232) <= not((inputs(212)) xor (inputs(75)));
    layer0_outputs(233) <= inputs(142);
    layer0_outputs(234) <= inputs(200);
    layer0_outputs(235) <= (inputs(132)) and not (inputs(78));
    layer0_outputs(236) <= inputs(131);
    layer0_outputs(237) <= not(inputs(120)) or (inputs(189));
    layer0_outputs(238) <= (inputs(189)) or (inputs(32));
    layer0_outputs(239) <= inputs(150);
    layer0_outputs(240) <= '0';
    layer0_outputs(241) <= inputs(245);
    layer0_outputs(242) <= (inputs(225)) or (inputs(150));
    layer0_outputs(243) <= inputs(127);
    layer0_outputs(244) <= '0';
    layer0_outputs(245) <= (inputs(133)) xor (inputs(186));
    layer0_outputs(246) <= not((inputs(171)) or (inputs(239)));
    layer0_outputs(247) <= (inputs(107)) and not (inputs(252));
    layer0_outputs(248) <= (inputs(185)) and not (inputs(208));
    layer0_outputs(249) <= (inputs(140)) xor (inputs(33));
    layer0_outputs(250) <= not((inputs(227)) or (inputs(193)));
    layer0_outputs(251) <= '1';
    layer0_outputs(252) <= not(inputs(172)) or (inputs(50));
    layer0_outputs(253) <= (inputs(146)) and (inputs(238));
    layer0_outputs(254) <= inputs(1);
    layer0_outputs(255) <= not(inputs(74)) or (inputs(78));
    layer0_outputs(256) <= inputs(124);
    layer0_outputs(257) <= inputs(152);
    layer0_outputs(258) <= (inputs(106)) and not (inputs(28));
    layer0_outputs(259) <= not(inputs(154));
    layer0_outputs(260) <= (inputs(219)) xor (inputs(160));
    layer0_outputs(261) <= not(inputs(87)) or (inputs(146));
    layer0_outputs(262) <= not(inputs(215)) or (inputs(41));
    layer0_outputs(263) <= (inputs(26)) xor (inputs(247));
    layer0_outputs(264) <= not(inputs(159));
    layer0_outputs(265) <= (inputs(200)) xor (inputs(63));
    layer0_outputs(266) <= inputs(68);
    layer0_outputs(267) <= not((inputs(138)) xor (inputs(223)));
    layer0_outputs(268) <= inputs(30);
    layer0_outputs(269) <= '0';
    layer0_outputs(270) <= not(inputs(120));
    layer0_outputs(271) <= (inputs(205)) xor (inputs(126));
    layer0_outputs(272) <= (inputs(230)) xor (inputs(36));
    layer0_outputs(273) <= (inputs(137)) and not (inputs(9));
    layer0_outputs(274) <= (inputs(72)) or (inputs(193));
    layer0_outputs(275) <= (inputs(68)) and not (inputs(221));
    layer0_outputs(276) <= not(inputs(92));
    layer0_outputs(277) <= (inputs(169)) and not (inputs(112));
    layer0_outputs(278) <= not((inputs(146)) or (inputs(82)));
    layer0_outputs(279) <= not((inputs(6)) and (inputs(17)));
    layer0_outputs(280) <= not(inputs(230));
    layer0_outputs(281) <= (inputs(115)) or (inputs(50));
    layer0_outputs(282) <= (inputs(92)) or (inputs(69));
    layer0_outputs(283) <= inputs(168);
    layer0_outputs(284) <= not((inputs(129)) and (inputs(31)));
    layer0_outputs(285) <= (inputs(236)) xor (inputs(0));
    layer0_outputs(286) <= not(inputs(254));
    layer0_outputs(287) <= (inputs(28)) or (inputs(163));
    layer0_outputs(288) <= not(inputs(122)) or (inputs(227));
    layer0_outputs(289) <= '1';
    layer0_outputs(290) <= not((inputs(155)) or (inputs(108)));
    layer0_outputs(291) <= not(inputs(167)) or (inputs(47));
    layer0_outputs(292) <= not((inputs(72)) or (inputs(98)));
    layer0_outputs(293) <= (inputs(179)) and not (inputs(22));
    layer0_outputs(294) <= '1';
    layer0_outputs(295) <= '0';
    layer0_outputs(296) <= (inputs(162)) and not (inputs(247));
    layer0_outputs(297) <= (inputs(135)) and not (inputs(33));
    layer0_outputs(298) <= (inputs(13)) or (inputs(165));
    layer0_outputs(299) <= (inputs(126)) and (inputs(115));
    layer0_outputs(300) <= not((inputs(82)) and (inputs(11)));
    layer0_outputs(301) <= (inputs(129)) xor (inputs(65));
    layer0_outputs(302) <= not(inputs(54)) or (inputs(133));
    layer0_outputs(303) <= not((inputs(37)) or (inputs(133)));
    layer0_outputs(304) <= not((inputs(23)) or (inputs(9)));
    layer0_outputs(305) <= (inputs(166)) and not (inputs(175));
    layer0_outputs(306) <= inputs(166);
    layer0_outputs(307) <= inputs(135);
    layer0_outputs(308) <= (inputs(8)) or (inputs(107));
    layer0_outputs(309) <= (inputs(137)) or (inputs(131));
    layer0_outputs(310) <= inputs(22);
    layer0_outputs(311) <= not(inputs(170));
    layer0_outputs(312) <= not(inputs(155));
    layer0_outputs(313) <= not(inputs(155));
    layer0_outputs(314) <= inputs(136);
    layer0_outputs(315) <= not(inputs(230)) or (inputs(1));
    layer0_outputs(316) <= inputs(120);
    layer0_outputs(317) <= not(inputs(168)) or (inputs(180));
    layer0_outputs(318) <= (inputs(192)) xor (inputs(191));
    layer0_outputs(319) <= not(inputs(87)) or (inputs(23));
    layer0_outputs(320) <= (inputs(170)) and not (inputs(51));
    layer0_outputs(321) <= (inputs(193)) xor (inputs(20));
    layer0_outputs(322) <= inputs(163);
    layer0_outputs(323) <= (inputs(106)) or (inputs(115));
    layer0_outputs(324) <= (inputs(220)) and (inputs(250));
    layer0_outputs(325) <= not(inputs(223));
    layer0_outputs(326) <= (inputs(58)) and not (inputs(104));
    layer0_outputs(327) <= (inputs(99)) or (inputs(98));
    layer0_outputs(328) <= not(inputs(106)) or (inputs(189));
    layer0_outputs(329) <= not(inputs(200));
    layer0_outputs(330) <= not(inputs(149)) or (inputs(129));
    layer0_outputs(331) <= (inputs(194)) xor (inputs(219));
    layer0_outputs(332) <= inputs(136);
    layer0_outputs(333) <= not((inputs(160)) and (inputs(254)));
    layer0_outputs(334) <= inputs(168);
    layer0_outputs(335) <= (inputs(165)) and not (inputs(14));
    layer0_outputs(336) <= not(inputs(184));
    layer0_outputs(337) <= not(inputs(215)) or (inputs(222));
    layer0_outputs(338) <= inputs(101);
    layer0_outputs(339) <= (inputs(90)) and not (inputs(108));
    layer0_outputs(340) <= not((inputs(185)) xor (inputs(15)));
    layer0_outputs(341) <= (inputs(214)) or (inputs(118));
    layer0_outputs(342) <= not(inputs(137)) or (inputs(4));
    layer0_outputs(343) <= inputs(71);
    layer0_outputs(344) <= inputs(33);
    layer0_outputs(345) <= not(inputs(133));
    layer0_outputs(346) <= inputs(177);
    layer0_outputs(347) <= (inputs(161)) or (inputs(163));
    layer0_outputs(348) <= not(inputs(131));
    layer0_outputs(349) <= not((inputs(161)) or (inputs(196)));
    layer0_outputs(350) <= inputs(181);
    layer0_outputs(351) <= not(inputs(246));
    layer0_outputs(352) <= not((inputs(158)) or (inputs(137)));
    layer0_outputs(353) <= not(inputs(196)) or (inputs(78));
    layer0_outputs(354) <= (inputs(4)) or (inputs(236));
    layer0_outputs(355) <= (inputs(209)) and not (inputs(160));
    layer0_outputs(356) <= (inputs(62)) or (inputs(76));
    layer0_outputs(357) <= (inputs(163)) and not (inputs(65));
    layer0_outputs(358) <= not((inputs(198)) or (inputs(167)));
    layer0_outputs(359) <= inputs(88);
    layer0_outputs(360) <= (inputs(152)) or (inputs(142));
    layer0_outputs(361) <= not((inputs(15)) xor (inputs(144)));
    layer0_outputs(362) <= (inputs(102)) or (inputs(12));
    layer0_outputs(363) <= not((inputs(147)) or (inputs(45)));
    layer0_outputs(364) <= (inputs(139)) or (inputs(112));
    layer0_outputs(365) <= inputs(171);
    layer0_outputs(366) <= not((inputs(69)) and (inputs(218)));
    layer0_outputs(367) <= (inputs(110)) or (inputs(102));
    layer0_outputs(368) <= not(inputs(178)) or (inputs(161));
    layer0_outputs(369) <= not(inputs(62)) or (inputs(11));
    layer0_outputs(370) <= not(inputs(152)) or (inputs(22));
    layer0_outputs(371) <= (inputs(115)) or (inputs(89));
    layer0_outputs(372) <= inputs(18);
    layer0_outputs(373) <= (inputs(121)) and not (inputs(40));
    layer0_outputs(374) <= (inputs(19)) and (inputs(33));
    layer0_outputs(375) <= (inputs(37)) or (inputs(24));
    layer0_outputs(376) <= not(inputs(214)) or (inputs(140));
    layer0_outputs(377) <= inputs(23);
    layer0_outputs(378) <= (inputs(220)) xor (inputs(50));
    layer0_outputs(379) <= (inputs(24)) xor (inputs(49));
    layer0_outputs(380) <= not((inputs(74)) xor (inputs(249)));
    layer0_outputs(381) <= not(inputs(30)) or (inputs(249));
    layer0_outputs(382) <= not(inputs(181));
    layer0_outputs(383) <= not(inputs(140));
    layer0_outputs(384) <= (inputs(174)) and not (inputs(48));
    layer0_outputs(385) <= not(inputs(150)) or (inputs(235));
    layer0_outputs(386) <= (inputs(147)) or (inputs(125));
    layer0_outputs(387) <= not(inputs(183));
    layer0_outputs(388) <= inputs(145);
    layer0_outputs(389) <= (inputs(188)) or (inputs(109));
    layer0_outputs(390) <= not(inputs(219));
    layer0_outputs(391) <= not(inputs(247)) or (inputs(1));
    layer0_outputs(392) <= not((inputs(178)) or (inputs(74)));
    layer0_outputs(393) <= '0';
    layer0_outputs(394) <= not(inputs(134));
    layer0_outputs(395) <= not((inputs(150)) or (inputs(108)));
    layer0_outputs(396) <= (inputs(145)) xor (inputs(232));
    layer0_outputs(397) <= not(inputs(153)) or (inputs(118));
    layer0_outputs(398) <= not((inputs(63)) xor (inputs(201)));
    layer0_outputs(399) <= (inputs(217)) or (inputs(171));
    layer0_outputs(400) <= (inputs(236)) xor (inputs(122));
    layer0_outputs(401) <= not(inputs(156));
    layer0_outputs(402) <= not((inputs(61)) xor (inputs(105)));
    layer0_outputs(403) <= inputs(139);
    layer0_outputs(404) <= (inputs(229)) xor (inputs(232));
    layer0_outputs(405) <= (inputs(237)) xor (inputs(27));
    layer0_outputs(406) <= not(inputs(196));
    layer0_outputs(407) <= (inputs(203)) and not (inputs(205));
    layer0_outputs(408) <= not(inputs(57));
    layer0_outputs(409) <= not((inputs(91)) or (inputs(81)));
    layer0_outputs(410) <= (inputs(219)) xor (inputs(222));
    layer0_outputs(411) <= inputs(124);
    layer0_outputs(412) <= inputs(147);
    layer0_outputs(413) <= not(inputs(118));
    layer0_outputs(414) <= not(inputs(86)) or (inputs(80));
    layer0_outputs(415) <= inputs(186);
    layer0_outputs(416) <= not((inputs(64)) and (inputs(204)));
    layer0_outputs(417) <= (inputs(253)) or (inputs(30));
    layer0_outputs(418) <= (inputs(244)) or (inputs(201));
    layer0_outputs(419) <= not(inputs(125));
    layer0_outputs(420) <= not(inputs(94)) or (inputs(13));
    layer0_outputs(421) <= not(inputs(75)) or (inputs(2));
    layer0_outputs(422) <= (inputs(231)) or (inputs(222));
    layer0_outputs(423) <= not(inputs(140));
    layer0_outputs(424) <= not((inputs(38)) or (inputs(195)));
    layer0_outputs(425) <= (inputs(107)) or (inputs(235));
    layer0_outputs(426) <= inputs(226);
    layer0_outputs(427) <= not(inputs(102)) or (inputs(80));
    layer0_outputs(428) <= not(inputs(135)) or (inputs(53));
    layer0_outputs(429) <= inputs(200);
    layer0_outputs(430) <= not(inputs(181));
    layer0_outputs(431) <= (inputs(63)) or (inputs(182));
    layer0_outputs(432) <= not(inputs(132));
    layer0_outputs(433) <= not((inputs(77)) or (inputs(250)));
    layer0_outputs(434) <= not(inputs(121)) or (inputs(24));
    layer0_outputs(435) <= not(inputs(24)) or (inputs(79));
    layer0_outputs(436) <= (inputs(144)) or (inputs(228));
    layer0_outputs(437) <= inputs(93);
    layer0_outputs(438) <= not((inputs(163)) or (inputs(39)));
    layer0_outputs(439) <= not((inputs(248)) or (inputs(124)));
    layer0_outputs(440) <= (inputs(119)) and not (inputs(146));
    layer0_outputs(441) <= not((inputs(128)) or (inputs(44)));
    layer0_outputs(442) <= '0';
    layer0_outputs(443) <= not(inputs(225));
    layer0_outputs(444) <= not(inputs(71)) or (inputs(205));
    layer0_outputs(445) <= not(inputs(23)) or (inputs(59));
    layer0_outputs(446) <= (inputs(122)) and not (inputs(250));
    layer0_outputs(447) <= not(inputs(58));
    layer0_outputs(448) <= not(inputs(141));
    layer0_outputs(449) <= not((inputs(70)) xor (inputs(222)));
    layer0_outputs(450) <= inputs(115);
    layer0_outputs(451) <= inputs(20);
    layer0_outputs(452) <= (inputs(219)) and not (inputs(2));
    layer0_outputs(453) <= (inputs(102)) xor (inputs(85));
    layer0_outputs(454) <= not((inputs(60)) xor (inputs(49)));
    layer0_outputs(455) <= (inputs(55)) or (inputs(141));
    layer0_outputs(456) <= (inputs(178)) or (inputs(39));
    layer0_outputs(457) <= not((inputs(51)) xor (inputs(28)));
    layer0_outputs(458) <= (inputs(179)) or (inputs(180));
    layer0_outputs(459) <= (inputs(94)) and not (inputs(11));
    layer0_outputs(460) <= inputs(77);
    layer0_outputs(461) <= (inputs(7)) and not (inputs(39));
    layer0_outputs(462) <= not((inputs(82)) or (inputs(253)));
    layer0_outputs(463) <= inputs(24);
    layer0_outputs(464) <= inputs(199);
    layer0_outputs(465) <= not(inputs(151));
    layer0_outputs(466) <= (inputs(103)) xor (inputs(64));
    layer0_outputs(467) <= not((inputs(116)) or (inputs(19)));
    layer0_outputs(468) <= (inputs(92)) and not (inputs(26));
    layer0_outputs(469) <= (inputs(151)) or (inputs(139));
    layer0_outputs(470) <= not(inputs(135));
    layer0_outputs(471) <= '0';
    layer0_outputs(472) <= inputs(185);
    layer0_outputs(473) <= not((inputs(188)) or (inputs(15)));
    layer0_outputs(474) <= not((inputs(125)) or (inputs(66)));
    layer0_outputs(475) <= '0';
    layer0_outputs(476) <= not(inputs(134)) or (inputs(149));
    layer0_outputs(477) <= not((inputs(127)) xor (inputs(177)));
    layer0_outputs(478) <= (inputs(79)) and not (inputs(142));
    layer0_outputs(479) <= not((inputs(37)) xor (inputs(243)));
    layer0_outputs(480) <= '0';
    layer0_outputs(481) <= inputs(94);
    layer0_outputs(482) <= (inputs(67)) xor (inputs(40));
    layer0_outputs(483) <= inputs(26);
    layer0_outputs(484) <= (inputs(90)) or (inputs(73));
    layer0_outputs(485) <= not((inputs(252)) or (inputs(167)));
    layer0_outputs(486) <= (inputs(158)) or (inputs(77));
    layer0_outputs(487) <= not((inputs(153)) or (inputs(53)));
    layer0_outputs(488) <= (inputs(60)) and not (inputs(234));
    layer0_outputs(489) <= not((inputs(26)) or (inputs(133)));
    layer0_outputs(490) <= (inputs(133)) and not (inputs(237));
    layer0_outputs(491) <= (inputs(77)) or (inputs(147));
    layer0_outputs(492) <= inputs(135);
    layer0_outputs(493) <= not(inputs(167));
    layer0_outputs(494) <= not(inputs(104)) or (inputs(171));
    layer0_outputs(495) <= (inputs(141)) and not (inputs(114));
    layer0_outputs(496) <= (inputs(141)) or (inputs(125));
    layer0_outputs(497) <= not(inputs(83));
    layer0_outputs(498) <= (inputs(85)) or (inputs(247));
    layer0_outputs(499) <= inputs(72);
    layer0_outputs(500) <= '0';
    layer0_outputs(501) <= '0';
    layer0_outputs(502) <= not((inputs(58)) xor (inputs(90)));
    layer0_outputs(503) <= not((inputs(26)) xor (inputs(251)));
    layer0_outputs(504) <= (inputs(255)) and not (inputs(175));
    layer0_outputs(505) <= not(inputs(247));
    layer0_outputs(506) <= (inputs(58)) xor (inputs(199));
    layer0_outputs(507) <= inputs(186);
    layer0_outputs(508) <= inputs(214);
    layer0_outputs(509) <= not(inputs(107));
    layer0_outputs(510) <= not(inputs(122));
    layer0_outputs(511) <= (inputs(58)) or (inputs(93));
    layer0_outputs(512) <= (inputs(159)) or (inputs(152));
    layer0_outputs(513) <= inputs(29);
    layer0_outputs(514) <= not(inputs(181)) or (inputs(177));
    layer0_outputs(515) <= (inputs(174)) xor (inputs(22));
    layer0_outputs(516) <= not((inputs(26)) or (inputs(164)));
    layer0_outputs(517) <= not((inputs(204)) xor (inputs(187)));
    layer0_outputs(518) <= '0';
    layer0_outputs(519) <= not(inputs(49)) or (inputs(128));
    layer0_outputs(520) <= (inputs(244)) xor (inputs(162));
    layer0_outputs(521) <= not((inputs(175)) xor (inputs(153)));
    layer0_outputs(522) <= inputs(150);
    layer0_outputs(523) <= (inputs(241)) xor (inputs(130));
    layer0_outputs(524) <= inputs(230);
    layer0_outputs(525) <= not(inputs(149)) or (inputs(163));
    layer0_outputs(526) <= '0';
    layer0_outputs(527) <= inputs(159);
    layer0_outputs(528) <= '0';
    layer0_outputs(529) <= not(inputs(165));
    layer0_outputs(530) <= not((inputs(205)) and (inputs(142)));
    layer0_outputs(531) <= not(inputs(100)) or (inputs(161));
    layer0_outputs(532) <= not(inputs(150)) or (inputs(25));
    layer0_outputs(533) <= not((inputs(103)) or (inputs(18)));
    layer0_outputs(534) <= not((inputs(153)) or (inputs(146)));
    layer0_outputs(535) <= not((inputs(163)) or (inputs(86)));
    layer0_outputs(536) <= not((inputs(253)) or (inputs(65)));
    layer0_outputs(537) <= (inputs(87)) or (inputs(179));
    layer0_outputs(538) <= not((inputs(57)) or (inputs(178)));
    layer0_outputs(539) <= (inputs(111)) and not (inputs(143));
    layer0_outputs(540) <= not((inputs(182)) or (inputs(148)));
    layer0_outputs(541) <= not((inputs(22)) or (inputs(121)));
    layer0_outputs(542) <= not(inputs(142)) or (inputs(80));
    layer0_outputs(543) <= not(inputs(185)) or (inputs(145));
    layer0_outputs(544) <= (inputs(97)) or (inputs(15));
    layer0_outputs(545) <= (inputs(37)) xor (inputs(113));
    layer0_outputs(546) <= (inputs(67)) or (inputs(54));
    layer0_outputs(547) <= not((inputs(235)) or (inputs(229)));
    layer0_outputs(548) <= not(inputs(200)) or (inputs(19));
    layer0_outputs(549) <= not(inputs(184)) or (inputs(255));
    layer0_outputs(550) <= not(inputs(186)) or (inputs(69));
    layer0_outputs(551) <= (inputs(212)) or (inputs(96));
    layer0_outputs(552) <= not(inputs(45)) or (inputs(160));
    layer0_outputs(553) <= (inputs(158)) or (inputs(27));
    layer0_outputs(554) <= not((inputs(223)) or (inputs(168)));
    layer0_outputs(555) <= (inputs(104)) and not (inputs(51));
    layer0_outputs(556) <= not(inputs(238)) or (inputs(158));
    layer0_outputs(557) <= not(inputs(156));
    layer0_outputs(558) <= not(inputs(164));
    layer0_outputs(559) <= '0';
    layer0_outputs(560) <= (inputs(104)) or (inputs(222));
    layer0_outputs(561) <= (inputs(71)) and not (inputs(82));
    layer0_outputs(562) <= not((inputs(153)) or (inputs(27)));
    layer0_outputs(563) <= not(inputs(7));
    layer0_outputs(564) <= '1';
    layer0_outputs(565) <= (inputs(22)) or (inputs(150));
    layer0_outputs(566) <= not(inputs(164)) or (inputs(130));
    layer0_outputs(567) <= not((inputs(147)) xor (inputs(192)));
    layer0_outputs(568) <= not((inputs(38)) or (inputs(197)));
    layer0_outputs(569) <= (inputs(145)) and not (inputs(176));
    layer0_outputs(570) <= inputs(40);
    layer0_outputs(571) <= not((inputs(3)) xor (inputs(228)));
    layer0_outputs(572) <= (inputs(237)) or (inputs(101));
    layer0_outputs(573) <= not(inputs(120));
    layer0_outputs(574) <= (inputs(114)) and (inputs(14));
    layer0_outputs(575) <= not(inputs(43)) or (inputs(174));
    layer0_outputs(576) <= (inputs(36)) and not (inputs(66));
    layer0_outputs(577) <= not(inputs(138));
    layer0_outputs(578) <= not(inputs(57)) or (inputs(162));
    layer0_outputs(579) <= not((inputs(145)) and (inputs(19)));
    layer0_outputs(580) <= inputs(131);
    layer0_outputs(581) <= (inputs(247)) or (inputs(98));
    layer0_outputs(582) <= (inputs(178)) or (inputs(78));
    layer0_outputs(583) <= (inputs(86)) and not (inputs(106));
    layer0_outputs(584) <= not(inputs(114)) or (inputs(191));
    layer0_outputs(585) <= (inputs(234)) and not (inputs(199));
    layer0_outputs(586) <= not((inputs(100)) or (inputs(115)));
    layer0_outputs(587) <= (inputs(226)) and not (inputs(14));
    layer0_outputs(588) <= '0';
    layer0_outputs(589) <= inputs(42);
    layer0_outputs(590) <= (inputs(95)) and (inputs(110));
    layer0_outputs(591) <= (inputs(112)) and not (inputs(227));
    layer0_outputs(592) <= '1';
    layer0_outputs(593) <= (inputs(153)) and not (inputs(13));
    layer0_outputs(594) <= not(inputs(88)) or (inputs(157));
    layer0_outputs(595) <= (inputs(10)) and not (inputs(95));
    layer0_outputs(596) <= not((inputs(35)) or (inputs(17)));
    layer0_outputs(597) <= not(inputs(17));
    layer0_outputs(598) <= (inputs(219)) xor (inputs(22));
    layer0_outputs(599) <= not(inputs(15));
    layer0_outputs(600) <= inputs(107);
    layer0_outputs(601) <= not(inputs(124)) or (inputs(237));
    layer0_outputs(602) <= not(inputs(168)) or (inputs(102));
    layer0_outputs(603) <= not((inputs(79)) and (inputs(174)));
    layer0_outputs(604) <= (inputs(211)) and not (inputs(2));
    layer0_outputs(605) <= inputs(98);
    layer0_outputs(606) <= (inputs(193)) and not (inputs(190));
    layer0_outputs(607) <= (inputs(35)) or (inputs(204));
    layer0_outputs(608) <= not((inputs(120)) xor (inputs(123)));
    layer0_outputs(609) <= (inputs(91)) or (inputs(240));
    layer0_outputs(610) <= not((inputs(192)) or (inputs(186)));
    layer0_outputs(611) <= (inputs(81)) and not (inputs(253));
    layer0_outputs(612) <= (inputs(119)) or (inputs(7));
    layer0_outputs(613) <= not(inputs(233)) or (inputs(34));
    layer0_outputs(614) <= (inputs(217)) or (inputs(93));
    layer0_outputs(615) <= not(inputs(248));
    layer0_outputs(616) <= not(inputs(123)) or (inputs(210));
    layer0_outputs(617) <= (inputs(227)) xor (inputs(212));
    layer0_outputs(618) <= not((inputs(46)) xor (inputs(35)));
    layer0_outputs(619) <= (inputs(179)) or (inputs(236));
    layer0_outputs(620) <= not((inputs(154)) or (inputs(179)));
    layer0_outputs(621) <= not(inputs(202)) or (inputs(189));
    layer0_outputs(622) <= (inputs(36)) or (inputs(96));
    layer0_outputs(623) <= (inputs(114)) and not (inputs(111));
    layer0_outputs(624) <= not(inputs(61));
    layer0_outputs(625) <= (inputs(91)) and not (inputs(248));
    layer0_outputs(626) <= inputs(103);
    layer0_outputs(627) <= inputs(186);
    layer0_outputs(628) <= (inputs(113)) xor (inputs(231));
    layer0_outputs(629) <= not(inputs(18)) or (inputs(248));
    layer0_outputs(630) <= inputs(104);
    layer0_outputs(631) <= not(inputs(25));
    layer0_outputs(632) <= (inputs(93)) and not (inputs(246));
    layer0_outputs(633) <= (inputs(50)) and not (inputs(130));
    layer0_outputs(634) <= (inputs(132)) and not (inputs(143));
    layer0_outputs(635) <= '1';
    layer0_outputs(636) <= not(inputs(62)) or (inputs(64));
    layer0_outputs(637) <= (inputs(230)) xor (inputs(178));
    layer0_outputs(638) <= not(inputs(184));
    layer0_outputs(639) <= not((inputs(69)) or (inputs(47)));
    layer0_outputs(640) <= not(inputs(84));
    layer0_outputs(641) <= (inputs(29)) xor (inputs(156));
    layer0_outputs(642) <= not((inputs(146)) or (inputs(130)));
    layer0_outputs(643) <= inputs(10);
    layer0_outputs(644) <= (inputs(46)) or (inputs(120));
    layer0_outputs(645) <= inputs(103);
    layer0_outputs(646) <= not((inputs(65)) xor (inputs(214)));
    layer0_outputs(647) <= (inputs(255)) and not (inputs(97));
    layer0_outputs(648) <= not(inputs(4));
    layer0_outputs(649) <= inputs(37);
    layer0_outputs(650) <= not((inputs(33)) or (inputs(33)));
    layer0_outputs(651) <= not(inputs(201)) or (inputs(146));
    layer0_outputs(652) <= (inputs(201)) and not (inputs(93));
    layer0_outputs(653) <= not((inputs(197)) xor (inputs(29)));
    layer0_outputs(654) <= inputs(60);
    layer0_outputs(655) <= not(inputs(105));
    layer0_outputs(656) <= not((inputs(82)) or (inputs(67)));
    layer0_outputs(657) <= '1';
    layer0_outputs(658) <= (inputs(17)) or (inputs(1));
    layer0_outputs(659) <= '0';
    layer0_outputs(660) <= (inputs(213)) and not (inputs(233));
    layer0_outputs(661) <= not(inputs(235));
    layer0_outputs(662) <= (inputs(52)) or (inputs(61));
    layer0_outputs(663) <= inputs(207);
    layer0_outputs(664) <= inputs(106);
    layer0_outputs(665) <= not((inputs(182)) xor (inputs(97)));
    layer0_outputs(666) <= inputs(85);
    layer0_outputs(667) <= not(inputs(172)) or (inputs(138));
    layer0_outputs(668) <= (inputs(12)) xor (inputs(187));
    layer0_outputs(669) <= not((inputs(141)) or (inputs(213)));
    layer0_outputs(670) <= not((inputs(51)) or (inputs(68)));
    layer0_outputs(671) <= (inputs(132)) and not (inputs(207));
    layer0_outputs(672) <= (inputs(149)) and not (inputs(5));
    layer0_outputs(673) <= not(inputs(209)) or (inputs(82));
    layer0_outputs(674) <= inputs(14);
    layer0_outputs(675) <= not((inputs(193)) and (inputs(67)));
    layer0_outputs(676) <= inputs(101);
    layer0_outputs(677) <= not((inputs(120)) xor (inputs(32)));
    layer0_outputs(678) <= not(inputs(183));
    layer0_outputs(679) <= '1';
    layer0_outputs(680) <= inputs(192);
    layer0_outputs(681) <= (inputs(68)) and not (inputs(24));
    layer0_outputs(682) <= (inputs(47)) xor (inputs(165));
    layer0_outputs(683) <= not((inputs(183)) xor (inputs(2)));
    layer0_outputs(684) <= not((inputs(195)) and (inputs(3)));
    layer0_outputs(685) <= '1';
    layer0_outputs(686) <= not(inputs(87));
    layer0_outputs(687) <= not(inputs(137)) or (inputs(57));
    layer0_outputs(688) <= not(inputs(151));
    layer0_outputs(689) <= not(inputs(121));
    layer0_outputs(690) <= not(inputs(239));
    layer0_outputs(691) <= inputs(117);
    layer0_outputs(692) <= inputs(218);
    layer0_outputs(693) <= (inputs(172)) and not (inputs(250));
    layer0_outputs(694) <= (inputs(110)) xor (inputs(203));
    layer0_outputs(695) <= not(inputs(11)) or (inputs(154));
    layer0_outputs(696) <= not(inputs(233)) or (inputs(15));
    layer0_outputs(697) <= (inputs(206)) and not (inputs(159));
    layer0_outputs(698) <= not(inputs(171)) or (inputs(244));
    layer0_outputs(699) <= not(inputs(6));
    layer0_outputs(700) <= (inputs(180)) and not (inputs(12));
    layer0_outputs(701) <= (inputs(194)) or (inputs(156));
    layer0_outputs(702) <= inputs(27);
    layer0_outputs(703) <= inputs(13);
    layer0_outputs(704) <= (inputs(41)) xor (inputs(39));
    layer0_outputs(705) <= not((inputs(93)) or (inputs(104)));
    layer0_outputs(706) <= (inputs(92)) and not (inputs(48));
    layer0_outputs(707) <= (inputs(169)) and not (inputs(128));
    layer0_outputs(708) <= '0';
    layer0_outputs(709) <= (inputs(249)) or (inputs(116));
    layer0_outputs(710) <= (inputs(228)) and not (inputs(2));
    layer0_outputs(711) <= (inputs(44)) and not (inputs(126));
    layer0_outputs(712) <= not((inputs(92)) or (inputs(214)));
    layer0_outputs(713) <= inputs(193);
    layer0_outputs(714) <= inputs(81);
    layer0_outputs(715) <= not(inputs(191));
    layer0_outputs(716) <= not(inputs(87));
    layer0_outputs(717) <= (inputs(5)) and (inputs(82));
    layer0_outputs(718) <= (inputs(191)) or (inputs(76));
    layer0_outputs(719) <= (inputs(110)) or (inputs(103));
    layer0_outputs(720) <= not((inputs(118)) or (inputs(139)));
    layer0_outputs(721) <= not(inputs(228));
    layer0_outputs(722) <= inputs(149);
    layer0_outputs(723) <= not((inputs(62)) or (inputs(170)));
    layer0_outputs(724) <= (inputs(233)) xor (inputs(25));
    layer0_outputs(725) <= (inputs(154)) or (inputs(173));
    layer0_outputs(726) <= not((inputs(52)) or (inputs(83)));
    layer0_outputs(727) <= '0';
    layer0_outputs(728) <= (inputs(85)) and not (inputs(51));
    layer0_outputs(729) <= (inputs(194)) or (inputs(40));
    layer0_outputs(730) <= (inputs(12)) xor (inputs(113));
    layer0_outputs(731) <= not((inputs(248)) and (inputs(236)));
    layer0_outputs(732) <= not(inputs(105));
    layer0_outputs(733) <= (inputs(86)) or (inputs(85));
    layer0_outputs(734) <= (inputs(199)) or (inputs(233));
    layer0_outputs(735) <= inputs(77);
    layer0_outputs(736) <= not(inputs(214));
    layer0_outputs(737) <= (inputs(117)) and not (inputs(246));
    layer0_outputs(738) <= (inputs(223)) xor (inputs(240));
    layer0_outputs(739) <= (inputs(94)) xor (inputs(186));
    layer0_outputs(740) <= not((inputs(219)) xor (inputs(53)));
    layer0_outputs(741) <= not(inputs(229));
    layer0_outputs(742) <= not(inputs(198)) or (inputs(209));
    layer0_outputs(743) <= (inputs(152)) and not (inputs(104));
    layer0_outputs(744) <= not((inputs(125)) or (inputs(196)));
    layer0_outputs(745) <= not(inputs(118));
    layer0_outputs(746) <= (inputs(155)) and not (inputs(49));
    layer0_outputs(747) <= not(inputs(155));
    layer0_outputs(748) <= not((inputs(96)) or (inputs(84)));
    layer0_outputs(749) <= not((inputs(114)) and (inputs(26)));
    layer0_outputs(750) <= not((inputs(53)) xor (inputs(127)));
    layer0_outputs(751) <= (inputs(117)) or (inputs(49));
    layer0_outputs(752) <= not(inputs(43)) or (inputs(5));
    layer0_outputs(753) <= (inputs(70)) and not (inputs(50));
    layer0_outputs(754) <= not((inputs(74)) and (inputs(200)));
    layer0_outputs(755) <= not((inputs(21)) or (inputs(234)));
    layer0_outputs(756) <= not((inputs(225)) or (inputs(13)));
    layer0_outputs(757) <= not(inputs(228)) or (inputs(19));
    layer0_outputs(758) <= (inputs(32)) xor (inputs(216));
    layer0_outputs(759) <= not(inputs(60));
    layer0_outputs(760) <= not((inputs(229)) or (inputs(39)));
    layer0_outputs(761) <= (inputs(37)) xor (inputs(82));
    layer0_outputs(762) <= not((inputs(37)) or (inputs(225)));
    layer0_outputs(763) <= (inputs(9)) xor (inputs(217));
    layer0_outputs(764) <= not((inputs(227)) or (inputs(136)));
    layer0_outputs(765) <= not((inputs(194)) or (inputs(111)));
    layer0_outputs(766) <= (inputs(241)) and (inputs(221));
    layer0_outputs(767) <= (inputs(26)) or (inputs(171));
    layer0_outputs(768) <= (inputs(24)) or (inputs(56));
    layer0_outputs(769) <= (inputs(201)) or (inputs(102));
    layer0_outputs(770) <= not(inputs(212)) or (inputs(135));
    layer0_outputs(771) <= inputs(63);
    layer0_outputs(772) <= inputs(82);
    layer0_outputs(773) <= not(inputs(123));
    layer0_outputs(774) <= inputs(32);
    layer0_outputs(775) <= (inputs(101)) and not (inputs(126));
    layer0_outputs(776) <= not((inputs(11)) xor (inputs(73)));
    layer0_outputs(777) <= (inputs(210)) and not (inputs(233));
    layer0_outputs(778) <= not((inputs(242)) or (inputs(41)));
    layer0_outputs(779) <= not(inputs(143));
    layer0_outputs(780) <= inputs(117);
    layer0_outputs(781) <= (inputs(193)) xor (inputs(243));
    layer0_outputs(782) <= (inputs(16)) xor (inputs(119));
    layer0_outputs(783) <= inputs(11);
    layer0_outputs(784) <= not(inputs(193)) or (inputs(81));
    layer0_outputs(785) <= not(inputs(89));
    layer0_outputs(786) <= '1';
    layer0_outputs(787) <= not((inputs(123)) or (inputs(132)));
    layer0_outputs(788) <= (inputs(2)) or (inputs(203));
    layer0_outputs(789) <= (inputs(160)) or (inputs(135));
    layer0_outputs(790) <= (inputs(198)) and (inputs(98));
    layer0_outputs(791) <= inputs(89);
    layer0_outputs(792) <= (inputs(66)) or (inputs(174));
    layer0_outputs(793) <= (inputs(115)) or (inputs(59));
    layer0_outputs(794) <= not((inputs(164)) or (inputs(136)));
    layer0_outputs(795) <= not(inputs(132));
    layer0_outputs(796) <= not((inputs(36)) xor (inputs(161)));
    layer0_outputs(797) <= not((inputs(52)) and (inputs(122)));
    layer0_outputs(798) <= not((inputs(237)) xor (inputs(157)));
    layer0_outputs(799) <= (inputs(40)) or (inputs(56));
    layer0_outputs(800) <= (inputs(58)) and not (inputs(6));
    layer0_outputs(801) <= not(inputs(73));
    layer0_outputs(802) <= (inputs(13)) or (inputs(175));
    layer0_outputs(803) <= not((inputs(180)) or (inputs(0)));
    layer0_outputs(804) <= not(inputs(137)) or (inputs(191));
    layer0_outputs(805) <= not((inputs(7)) or (inputs(201)));
    layer0_outputs(806) <= not(inputs(114)) or (inputs(21));
    layer0_outputs(807) <= inputs(32);
    layer0_outputs(808) <= (inputs(32)) and (inputs(15));
    layer0_outputs(809) <= not((inputs(25)) xor (inputs(104)));
    layer0_outputs(810) <= (inputs(170)) or (inputs(210));
    layer0_outputs(811) <= (inputs(146)) or (inputs(10));
    layer0_outputs(812) <= not((inputs(187)) xor (inputs(19)));
    layer0_outputs(813) <= not((inputs(71)) and (inputs(2)));
    layer0_outputs(814) <= not((inputs(29)) and (inputs(132)));
    layer0_outputs(815) <= (inputs(190)) xor (inputs(80));
    layer0_outputs(816) <= not((inputs(152)) xor (inputs(11)));
    layer0_outputs(817) <= (inputs(129)) xor (inputs(121));
    layer0_outputs(818) <= not((inputs(232)) xor (inputs(64)));
    layer0_outputs(819) <= '0';
    layer0_outputs(820) <= '1';
    layer0_outputs(821) <= not(inputs(122)) or (inputs(61));
    layer0_outputs(822) <= not(inputs(57));
    layer0_outputs(823) <= not((inputs(95)) xor (inputs(182)));
    layer0_outputs(824) <= not(inputs(83)) or (inputs(157));
    layer0_outputs(825) <= '1';
    layer0_outputs(826) <= inputs(67);
    layer0_outputs(827) <= (inputs(116)) or (inputs(135));
    layer0_outputs(828) <= not((inputs(108)) or (inputs(50)));
    layer0_outputs(829) <= not(inputs(155));
    layer0_outputs(830) <= not(inputs(100));
    layer0_outputs(831) <= not(inputs(122));
    layer0_outputs(832) <= not(inputs(48));
    layer0_outputs(833) <= not(inputs(254));
    layer0_outputs(834) <= (inputs(59)) and not (inputs(5));
    layer0_outputs(835) <= '0';
    layer0_outputs(836) <= not(inputs(205));
    layer0_outputs(837) <= not(inputs(217));
    layer0_outputs(838) <= not((inputs(171)) or (inputs(40)));
    layer0_outputs(839) <= not((inputs(47)) and (inputs(153)));
    layer0_outputs(840) <= not(inputs(102));
    layer0_outputs(841) <= not((inputs(199)) and (inputs(167)));
    layer0_outputs(842) <= not(inputs(228));
    layer0_outputs(843) <= (inputs(88)) or (inputs(23));
    layer0_outputs(844) <= not(inputs(152));
    layer0_outputs(845) <= (inputs(252)) and not (inputs(213));
    layer0_outputs(846) <= not((inputs(114)) and (inputs(103)));
    layer0_outputs(847) <= (inputs(81)) and not (inputs(255));
    layer0_outputs(848) <= (inputs(78)) or (inputs(234));
    layer0_outputs(849) <= not(inputs(27));
    layer0_outputs(850) <= not(inputs(131));
    layer0_outputs(851) <= not(inputs(60)) or (inputs(223));
    layer0_outputs(852) <= '1';
    layer0_outputs(853) <= not(inputs(119));
    layer0_outputs(854) <= '0';
    layer0_outputs(855) <= (inputs(134)) and not (inputs(59));
    layer0_outputs(856) <= (inputs(153)) or (inputs(83));
    layer0_outputs(857) <= not((inputs(203)) or (inputs(196)));
    layer0_outputs(858) <= (inputs(35)) and (inputs(207));
    layer0_outputs(859) <= not(inputs(32));
    layer0_outputs(860) <= not((inputs(101)) or (inputs(224)));
    layer0_outputs(861) <= not(inputs(92));
    layer0_outputs(862) <= (inputs(38)) and not (inputs(81));
    layer0_outputs(863) <= (inputs(167)) or (inputs(100));
    layer0_outputs(864) <= inputs(54);
    layer0_outputs(865) <= not(inputs(27));
    layer0_outputs(866) <= (inputs(254)) xor (inputs(86));
    layer0_outputs(867) <= (inputs(244)) and not (inputs(128));
    layer0_outputs(868) <= not((inputs(132)) and (inputs(10)));
    layer0_outputs(869) <= (inputs(113)) and not (inputs(237));
    layer0_outputs(870) <= not((inputs(154)) or (inputs(200)));
    layer0_outputs(871) <= not((inputs(172)) or (inputs(215)));
    layer0_outputs(872) <= not((inputs(140)) or (inputs(42)));
    layer0_outputs(873) <= not((inputs(21)) or (inputs(195)));
    layer0_outputs(874) <= not(inputs(153));
    layer0_outputs(875) <= (inputs(125)) and not (inputs(8));
    layer0_outputs(876) <= not((inputs(64)) and (inputs(222)));
    layer0_outputs(877) <= not((inputs(196)) or (inputs(82)));
    layer0_outputs(878) <= not(inputs(250));
    layer0_outputs(879) <= (inputs(139)) and not (inputs(45));
    layer0_outputs(880) <= not(inputs(72));
    layer0_outputs(881) <= (inputs(148)) and not (inputs(215));
    layer0_outputs(882) <= not(inputs(84)) or (inputs(159));
    layer0_outputs(883) <= not((inputs(157)) or (inputs(123)));
    layer0_outputs(884) <= inputs(138);
    layer0_outputs(885) <= not((inputs(201)) or (inputs(220)));
    layer0_outputs(886) <= not(inputs(171)) or (inputs(126));
    layer0_outputs(887) <= not(inputs(11)) or (inputs(124));
    layer0_outputs(888) <= (inputs(123)) or (inputs(221));
    layer0_outputs(889) <= (inputs(151)) and not (inputs(113));
    layer0_outputs(890) <= not((inputs(30)) xor (inputs(30)));
    layer0_outputs(891) <= not(inputs(38));
    layer0_outputs(892) <= not((inputs(173)) xor (inputs(247)));
    layer0_outputs(893) <= not(inputs(6)) or (inputs(10));
    layer0_outputs(894) <= (inputs(244)) xor (inputs(85));
    layer0_outputs(895) <= not((inputs(166)) or (inputs(82)));
    layer0_outputs(896) <= not(inputs(185)) or (inputs(93));
    layer0_outputs(897) <= not((inputs(249)) or (inputs(233)));
    layer0_outputs(898) <= not(inputs(234)) or (inputs(208));
    layer0_outputs(899) <= not(inputs(156));
    layer0_outputs(900) <= not((inputs(103)) or (inputs(186)));
    layer0_outputs(901) <= not(inputs(232)) or (inputs(173));
    layer0_outputs(902) <= not((inputs(95)) and (inputs(190)));
    layer0_outputs(903) <= not((inputs(180)) or (inputs(220)));
    layer0_outputs(904) <= not(inputs(149));
    layer0_outputs(905) <= not(inputs(98));
    layer0_outputs(906) <= (inputs(139)) and not (inputs(206));
    layer0_outputs(907) <= (inputs(85)) and not (inputs(187));
    layer0_outputs(908) <= not((inputs(151)) or (inputs(225)));
    layer0_outputs(909) <= not(inputs(42));
    layer0_outputs(910) <= not(inputs(85));
    layer0_outputs(911) <= not((inputs(189)) xor (inputs(143)));
    layer0_outputs(912) <= '0';
    layer0_outputs(913) <= '0';
    layer0_outputs(914) <= not(inputs(186)) or (inputs(128));
    layer0_outputs(915) <= not((inputs(90)) and (inputs(199)));
    layer0_outputs(916) <= inputs(122);
    layer0_outputs(917) <= (inputs(74)) and not (inputs(247));
    layer0_outputs(918) <= (inputs(17)) xor (inputs(211));
    layer0_outputs(919) <= inputs(116);
    layer0_outputs(920) <= inputs(43);
    layer0_outputs(921) <= not(inputs(149));
    layer0_outputs(922) <= (inputs(147)) or (inputs(61));
    layer0_outputs(923) <= not((inputs(164)) or (inputs(79)));
    layer0_outputs(924) <= inputs(90);
    layer0_outputs(925) <= not(inputs(177)) or (inputs(238));
    layer0_outputs(926) <= not((inputs(113)) xor (inputs(150)));
    layer0_outputs(927) <= not((inputs(125)) or (inputs(141)));
    layer0_outputs(928) <= (inputs(196)) and not (inputs(100));
    layer0_outputs(929) <= not((inputs(21)) or (inputs(105)));
    layer0_outputs(930) <= not(inputs(199)) or (inputs(130));
    layer0_outputs(931) <= not(inputs(25));
    layer0_outputs(932) <= not((inputs(124)) or (inputs(48)));
    layer0_outputs(933) <= (inputs(180)) and not (inputs(159));
    layer0_outputs(934) <= inputs(183);
    layer0_outputs(935) <= inputs(102);
    layer0_outputs(936) <= not(inputs(57));
    layer0_outputs(937) <= not(inputs(122)) or (inputs(202));
    layer0_outputs(938) <= (inputs(20)) xor (inputs(251));
    layer0_outputs(939) <= not(inputs(117));
    layer0_outputs(940) <= (inputs(165)) or (inputs(189));
    layer0_outputs(941) <= not(inputs(166));
    layer0_outputs(942) <= not(inputs(185));
    layer0_outputs(943) <= not(inputs(138)) or (inputs(193));
    layer0_outputs(944) <= (inputs(216)) and not (inputs(25));
    layer0_outputs(945) <= not(inputs(24));
    layer0_outputs(946) <= not((inputs(112)) xor (inputs(198)));
    layer0_outputs(947) <= inputs(235);
    layer0_outputs(948) <= not((inputs(106)) or (inputs(235)));
    layer0_outputs(949) <= not((inputs(194)) or (inputs(71)));
    layer0_outputs(950) <= '1';
    layer0_outputs(951) <= not((inputs(3)) and (inputs(228)));
    layer0_outputs(952) <= not((inputs(178)) or (inputs(89)));
    layer0_outputs(953) <= not((inputs(207)) and (inputs(236)));
    layer0_outputs(954) <= not(inputs(121));
    layer0_outputs(955) <= (inputs(189)) or (inputs(54));
    layer0_outputs(956) <= (inputs(21)) xor (inputs(190));
    layer0_outputs(957) <= not((inputs(47)) and (inputs(65)));
    layer0_outputs(958) <= inputs(182);
    layer0_outputs(959) <= not((inputs(194)) and (inputs(246)));
    layer0_outputs(960) <= not((inputs(130)) xor (inputs(84)));
    layer0_outputs(961) <= (inputs(74)) and not (inputs(255));
    layer0_outputs(962) <= (inputs(15)) xor (inputs(10));
    layer0_outputs(963) <= not(inputs(26));
    layer0_outputs(964) <= inputs(204);
    layer0_outputs(965) <= (inputs(51)) or (inputs(180));
    layer0_outputs(966) <= inputs(5);
    layer0_outputs(967) <= (inputs(49)) xor (inputs(66));
    layer0_outputs(968) <= not((inputs(114)) or (inputs(14)));
    layer0_outputs(969) <= not(inputs(181));
    layer0_outputs(970) <= (inputs(113)) and not (inputs(30));
    layer0_outputs(971) <= not(inputs(113));
    layer0_outputs(972) <= not((inputs(62)) xor (inputs(176)));
    layer0_outputs(973) <= not((inputs(216)) or (inputs(232)));
    layer0_outputs(974) <= not(inputs(248));
    layer0_outputs(975) <= (inputs(168)) or (inputs(7));
    layer0_outputs(976) <= inputs(86);
    layer0_outputs(977) <= inputs(44);
    layer0_outputs(978) <= (inputs(80)) and (inputs(212));
    layer0_outputs(979) <= not(inputs(192));
    layer0_outputs(980) <= not(inputs(196));
    layer0_outputs(981) <= (inputs(41)) and not (inputs(12));
    layer0_outputs(982) <= not(inputs(72));
    layer0_outputs(983) <= inputs(153);
    layer0_outputs(984) <= (inputs(254)) xor (inputs(40));
    layer0_outputs(985) <= not(inputs(76));
    layer0_outputs(986) <= (inputs(180)) or (inputs(157));
    layer0_outputs(987) <= not((inputs(147)) or (inputs(163)));
    layer0_outputs(988) <= not((inputs(33)) xor (inputs(224)));
    layer0_outputs(989) <= (inputs(56)) or (inputs(118));
    layer0_outputs(990) <= not((inputs(128)) and (inputs(80)));
    layer0_outputs(991) <= (inputs(153)) and not (inputs(212));
    layer0_outputs(992) <= not((inputs(111)) or (inputs(74)));
    layer0_outputs(993) <= not((inputs(186)) and (inputs(214)));
    layer0_outputs(994) <= '1';
    layer0_outputs(995) <= (inputs(200)) and not (inputs(206));
    layer0_outputs(996) <= not((inputs(203)) xor (inputs(114)));
    layer0_outputs(997) <= not(inputs(31)) or (inputs(37));
    layer0_outputs(998) <= inputs(104);
    layer0_outputs(999) <= (inputs(89)) or (inputs(162));
    layer0_outputs(1000) <= not((inputs(233)) or (inputs(182)));
    layer0_outputs(1001) <= (inputs(91)) or (inputs(80));
    layer0_outputs(1002) <= (inputs(78)) xor (inputs(2));
    layer0_outputs(1003) <= not((inputs(104)) or (inputs(48)));
    layer0_outputs(1004) <= (inputs(26)) or (inputs(38));
    layer0_outputs(1005) <= not((inputs(9)) or (inputs(36)));
    layer0_outputs(1006) <= not((inputs(148)) or (inputs(121)));
    layer0_outputs(1007) <= not(inputs(197));
    layer0_outputs(1008) <= not((inputs(247)) xor (inputs(229)));
    layer0_outputs(1009) <= not(inputs(230));
    layer0_outputs(1010) <= (inputs(134)) xor (inputs(9));
    layer0_outputs(1011) <= (inputs(190)) or (inputs(178));
    layer0_outputs(1012) <= not(inputs(56));
    layer0_outputs(1013) <= '1';
    layer0_outputs(1014) <= not(inputs(225)) or (inputs(120));
    layer0_outputs(1015) <= not(inputs(223));
    layer0_outputs(1016) <= inputs(27);
    layer0_outputs(1017) <= not(inputs(240));
    layer0_outputs(1018) <= not((inputs(14)) or (inputs(40)));
    layer0_outputs(1019) <= (inputs(68)) and not (inputs(11));
    layer0_outputs(1020) <= (inputs(51)) and (inputs(191));
    layer0_outputs(1021) <= not((inputs(251)) and (inputs(8)));
    layer0_outputs(1022) <= (inputs(83)) or (inputs(174));
    layer0_outputs(1023) <= not(inputs(199));
    layer0_outputs(1024) <= (inputs(123)) or (inputs(95));
    layer0_outputs(1025) <= '1';
    layer0_outputs(1026) <= (inputs(184)) xor (inputs(10));
    layer0_outputs(1027) <= inputs(14);
    layer0_outputs(1028) <= not((inputs(43)) or (inputs(139)));
    layer0_outputs(1029) <= '0';
    layer0_outputs(1030) <= inputs(141);
    layer0_outputs(1031) <= (inputs(93)) or (inputs(191));
    layer0_outputs(1032) <= '1';
    layer0_outputs(1033) <= (inputs(71)) and not (inputs(60));
    layer0_outputs(1034) <= not((inputs(76)) or (inputs(202)));
    layer0_outputs(1035) <= (inputs(202)) or (inputs(28));
    layer0_outputs(1036) <= not((inputs(59)) or (inputs(128)));
    layer0_outputs(1037) <= inputs(151);
    layer0_outputs(1038) <= (inputs(248)) or (inputs(228));
    layer0_outputs(1039) <= (inputs(12)) xor (inputs(203));
    layer0_outputs(1040) <= not((inputs(23)) or (inputs(230)));
    layer0_outputs(1041) <= not(inputs(134));
    layer0_outputs(1042) <= not((inputs(146)) or (inputs(134)));
    layer0_outputs(1043) <= not(inputs(183)) or (inputs(178));
    layer0_outputs(1044) <= (inputs(58)) and not (inputs(250));
    layer0_outputs(1045) <= (inputs(171)) xor (inputs(193));
    layer0_outputs(1046) <= not((inputs(190)) or (inputs(136)));
    layer0_outputs(1047) <= (inputs(96)) xor (inputs(225));
    layer0_outputs(1048) <= (inputs(140)) or (inputs(232));
    layer0_outputs(1049) <= (inputs(203)) or (inputs(196));
    layer0_outputs(1050) <= (inputs(126)) xor (inputs(89));
    layer0_outputs(1051) <= '0';
    layer0_outputs(1052) <= inputs(230);
    layer0_outputs(1053) <= (inputs(90)) and not (inputs(99));
    layer0_outputs(1054) <= '0';
    layer0_outputs(1055) <= not((inputs(64)) xor (inputs(226)));
    layer0_outputs(1056) <= (inputs(161)) or (inputs(106));
    layer0_outputs(1057) <= (inputs(89)) or (inputs(77));
    layer0_outputs(1058) <= not((inputs(161)) and (inputs(226)));
    layer0_outputs(1059) <= not((inputs(63)) xor (inputs(189)));
    layer0_outputs(1060) <= (inputs(109)) or (inputs(47));
    layer0_outputs(1061) <= (inputs(167)) and (inputs(137));
    layer0_outputs(1062) <= (inputs(200)) or (inputs(109));
    layer0_outputs(1063) <= not(inputs(94)) or (inputs(144));
    layer0_outputs(1064) <= (inputs(42)) and not (inputs(9));
    layer0_outputs(1065) <= '0';
    layer0_outputs(1066) <= (inputs(65)) or (inputs(162));
    layer0_outputs(1067) <= (inputs(138)) and not (inputs(234));
    layer0_outputs(1068) <= not(inputs(72)) or (inputs(224));
    layer0_outputs(1069) <= not(inputs(136)) or (inputs(23));
    layer0_outputs(1070) <= (inputs(179)) and not (inputs(66));
    layer0_outputs(1071) <= not(inputs(41));
    layer0_outputs(1072) <= '0';
    layer0_outputs(1073) <= not((inputs(234)) or (inputs(9)));
    layer0_outputs(1074) <= inputs(105);
    layer0_outputs(1075) <= not((inputs(41)) xor (inputs(156)));
    layer0_outputs(1076) <= (inputs(244)) xor (inputs(125));
    layer0_outputs(1077) <= not(inputs(251));
    layer0_outputs(1078) <= not((inputs(83)) or (inputs(97)));
    layer0_outputs(1079) <= not((inputs(189)) or (inputs(189)));
    layer0_outputs(1080) <= (inputs(195)) and not (inputs(223));
    layer0_outputs(1081) <= not((inputs(202)) xor (inputs(146)));
    layer0_outputs(1082) <= (inputs(57)) and not (inputs(63));
    layer0_outputs(1083) <= not(inputs(119)) or (inputs(142));
    layer0_outputs(1084) <= (inputs(36)) and not (inputs(95));
    layer0_outputs(1085) <= not(inputs(33)) or (inputs(112));
    layer0_outputs(1086) <= not((inputs(35)) or (inputs(122)));
    layer0_outputs(1087) <= not((inputs(92)) or (inputs(40)));
    layer0_outputs(1088) <= (inputs(113)) and (inputs(110));
    layer0_outputs(1089) <= (inputs(64)) and not (inputs(114));
    layer0_outputs(1090) <= (inputs(197)) and not (inputs(97));
    layer0_outputs(1091) <= not((inputs(64)) xor (inputs(141)));
    layer0_outputs(1092) <= (inputs(169)) and not (inputs(44));
    layer0_outputs(1093) <= (inputs(174)) and not (inputs(176));
    layer0_outputs(1094) <= inputs(99);
    layer0_outputs(1095) <= not(inputs(6)) or (inputs(143));
    layer0_outputs(1096) <= not(inputs(68));
    layer0_outputs(1097) <= not(inputs(176)) or (inputs(33));
    layer0_outputs(1098) <= not((inputs(140)) or (inputs(186)));
    layer0_outputs(1099) <= not((inputs(172)) or (inputs(155)));
    layer0_outputs(1100) <= not((inputs(66)) or (inputs(137)));
    layer0_outputs(1101) <= not((inputs(28)) xor (inputs(47)));
    layer0_outputs(1102) <= not(inputs(163));
    layer0_outputs(1103) <= (inputs(169)) and not (inputs(45));
    layer0_outputs(1104) <= inputs(89);
    layer0_outputs(1105) <= (inputs(205)) or (inputs(54));
    layer0_outputs(1106) <= not((inputs(30)) xor (inputs(60)));
    layer0_outputs(1107) <= (inputs(81)) xor (inputs(60));
    layer0_outputs(1108) <= not(inputs(39));
    layer0_outputs(1109) <= not(inputs(97)) or (inputs(62));
    layer0_outputs(1110) <= inputs(252);
    layer0_outputs(1111) <= (inputs(149)) and (inputs(185));
    layer0_outputs(1112) <= (inputs(170)) and (inputs(75));
    layer0_outputs(1113) <= not((inputs(232)) xor (inputs(240)));
    layer0_outputs(1114) <= not(inputs(173)) or (inputs(50));
    layer0_outputs(1115) <= not(inputs(148));
    layer0_outputs(1116) <= inputs(203);
    layer0_outputs(1117) <= not((inputs(255)) xor (inputs(165)));
    layer0_outputs(1118) <= (inputs(13)) and not (inputs(79));
    layer0_outputs(1119) <= inputs(105);
    layer0_outputs(1120) <= not(inputs(239)) or (inputs(214));
    layer0_outputs(1121) <= inputs(53);
    layer0_outputs(1122) <= (inputs(172)) and not (inputs(245));
    layer0_outputs(1123) <= '1';
    layer0_outputs(1124) <= not(inputs(108)) or (inputs(46));
    layer0_outputs(1125) <= inputs(234);
    layer0_outputs(1126) <= (inputs(42)) and not (inputs(195));
    layer0_outputs(1127) <= (inputs(161)) xor (inputs(240));
    layer0_outputs(1128) <= (inputs(75)) xor (inputs(177));
    layer0_outputs(1129) <= not(inputs(61)) or (inputs(23));
    layer0_outputs(1130) <= (inputs(85)) or (inputs(94));
    layer0_outputs(1131) <= (inputs(59)) and not (inputs(142));
    layer0_outputs(1132) <= (inputs(42)) xor (inputs(15));
    layer0_outputs(1133) <= inputs(200);
    layer0_outputs(1134) <= (inputs(215)) and not (inputs(66));
    layer0_outputs(1135) <= not(inputs(59));
    layer0_outputs(1136) <= not((inputs(82)) or (inputs(235)));
    layer0_outputs(1137) <= not((inputs(247)) and (inputs(250)));
    layer0_outputs(1138) <= (inputs(102)) and not (inputs(244));
    layer0_outputs(1139) <= (inputs(202)) xor (inputs(142));
    layer0_outputs(1140) <= inputs(177);
    layer0_outputs(1141) <= not(inputs(135)) or (inputs(253));
    layer0_outputs(1142) <= not((inputs(16)) or (inputs(109)));
    layer0_outputs(1143) <= not(inputs(37));
    layer0_outputs(1144) <= (inputs(127)) xor (inputs(215));
    layer0_outputs(1145) <= not(inputs(44)) or (inputs(192));
    layer0_outputs(1146) <= not((inputs(81)) or (inputs(50)));
    layer0_outputs(1147) <= inputs(17);
    layer0_outputs(1148) <= inputs(232);
    layer0_outputs(1149) <= (inputs(104)) and not (inputs(48));
    layer0_outputs(1150) <= not(inputs(100)) or (inputs(60));
    layer0_outputs(1151) <= not(inputs(44));
    layer0_outputs(1152) <= not(inputs(86)) or (inputs(158));
    layer0_outputs(1153) <= inputs(238);
    layer0_outputs(1154) <= not(inputs(58));
    layer0_outputs(1155) <= not(inputs(52));
    layer0_outputs(1156) <= not((inputs(211)) or (inputs(178)));
    layer0_outputs(1157) <= not((inputs(131)) or (inputs(245)));
    layer0_outputs(1158) <= inputs(232);
    layer0_outputs(1159) <= not(inputs(39)) or (inputs(62));
    layer0_outputs(1160) <= (inputs(136)) and not (inputs(28));
    layer0_outputs(1161) <= (inputs(60)) and (inputs(52));
    layer0_outputs(1162) <= '0';
    layer0_outputs(1163) <= (inputs(59)) xor (inputs(0));
    layer0_outputs(1164) <= not((inputs(116)) or (inputs(208)));
    layer0_outputs(1165) <= not(inputs(150));
    layer0_outputs(1166) <= (inputs(106)) and not (inputs(239));
    layer0_outputs(1167) <= not((inputs(36)) or (inputs(41)));
    layer0_outputs(1168) <= (inputs(58)) and not (inputs(241));
    layer0_outputs(1169) <= inputs(139);
    layer0_outputs(1170) <= (inputs(95)) xor (inputs(231));
    layer0_outputs(1171) <= (inputs(57)) or (inputs(203));
    layer0_outputs(1172) <= (inputs(46)) and not (inputs(63));
    layer0_outputs(1173) <= not(inputs(187));
    layer0_outputs(1174) <= (inputs(236)) and not (inputs(112));
    layer0_outputs(1175) <= (inputs(244)) and not (inputs(124));
    layer0_outputs(1176) <= inputs(114);
    layer0_outputs(1177) <= not((inputs(92)) xor (inputs(109)));
    layer0_outputs(1178) <= not((inputs(72)) or (inputs(113)));
    layer0_outputs(1179) <= inputs(175);
    layer0_outputs(1180) <= (inputs(47)) xor (inputs(125));
    layer0_outputs(1181) <= not((inputs(246)) or (inputs(158)));
    layer0_outputs(1182) <= not(inputs(213)) or (inputs(141));
    layer0_outputs(1183) <= '1';
    layer0_outputs(1184) <= (inputs(31)) xor (inputs(191));
    layer0_outputs(1185) <= not(inputs(6));
    layer0_outputs(1186) <= not(inputs(142)) or (inputs(59));
    layer0_outputs(1187) <= not((inputs(72)) or (inputs(234)));
    layer0_outputs(1188) <= (inputs(69)) xor (inputs(246));
    layer0_outputs(1189) <= not(inputs(194)) or (inputs(199));
    layer0_outputs(1190) <= (inputs(89)) and not (inputs(55));
    layer0_outputs(1191) <= not(inputs(239)) or (inputs(126));
    layer0_outputs(1192) <= inputs(86);
    layer0_outputs(1193) <= not(inputs(54)) or (inputs(113));
    layer0_outputs(1194) <= (inputs(243)) and (inputs(238));
    layer0_outputs(1195) <= (inputs(117)) xor (inputs(226));
    layer0_outputs(1196) <= (inputs(215)) or (inputs(55));
    layer0_outputs(1197) <= not(inputs(157));
    layer0_outputs(1198) <= not((inputs(240)) xor (inputs(21)));
    layer0_outputs(1199) <= not((inputs(215)) or (inputs(50)));
    layer0_outputs(1200) <= inputs(91);
    layer0_outputs(1201) <= not(inputs(200));
    layer0_outputs(1202) <= (inputs(52)) xor (inputs(76));
    layer0_outputs(1203) <= (inputs(172)) xor (inputs(80));
    layer0_outputs(1204) <= inputs(142);
    layer0_outputs(1205) <= inputs(108);
    layer0_outputs(1206) <= not(inputs(212));
    layer0_outputs(1207) <= inputs(205);
    layer0_outputs(1208) <= (inputs(252)) and not (inputs(43));
    layer0_outputs(1209) <= not(inputs(229));
    layer0_outputs(1210) <= not(inputs(153));
    layer0_outputs(1211) <= not(inputs(134)) or (inputs(104));
    layer0_outputs(1212) <= '0';
    layer0_outputs(1213) <= not((inputs(23)) or (inputs(141)));
    layer0_outputs(1214) <= inputs(141);
    layer0_outputs(1215) <= not(inputs(87));
    layer0_outputs(1216) <= not(inputs(182));
    layer0_outputs(1217) <= inputs(45);
    layer0_outputs(1218) <= '0';
    layer0_outputs(1219) <= not(inputs(73)) or (inputs(44));
    layer0_outputs(1220) <= inputs(241);
    layer0_outputs(1221) <= (inputs(18)) and (inputs(130));
    layer0_outputs(1222) <= not(inputs(70));
    layer0_outputs(1223) <= not(inputs(113));
    layer0_outputs(1224) <= (inputs(223)) and (inputs(52));
    layer0_outputs(1225) <= not(inputs(77)) or (inputs(239));
    layer0_outputs(1226) <= not((inputs(169)) or (inputs(205)));
    layer0_outputs(1227) <= not((inputs(151)) or (inputs(152)));
    layer0_outputs(1228) <= inputs(82);
    layer0_outputs(1229) <= not(inputs(54)) or (inputs(164));
    layer0_outputs(1230) <= not(inputs(132));
    layer0_outputs(1231) <= (inputs(70)) and not (inputs(68));
    layer0_outputs(1232) <= (inputs(67)) xor (inputs(226));
    layer0_outputs(1233) <= (inputs(173)) and not (inputs(110));
    layer0_outputs(1234) <= (inputs(66)) or (inputs(92));
    layer0_outputs(1235) <= '0';
    layer0_outputs(1236) <= not(inputs(170));
    layer0_outputs(1237) <= inputs(43);
    layer0_outputs(1238) <= (inputs(3)) or (inputs(149));
    layer0_outputs(1239) <= (inputs(13)) and not (inputs(219));
    layer0_outputs(1240) <= inputs(205);
    layer0_outputs(1241) <= not((inputs(188)) or (inputs(231)));
    layer0_outputs(1242) <= not(inputs(103)) or (inputs(193));
    layer0_outputs(1243) <= (inputs(129)) or (inputs(231));
    layer0_outputs(1244) <= inputs(182);
    layer0_outputs(1245) <= (inputs(133)) or (inputs(116));
    layer0_outputs(1246) <= '0';
    layer0_outputs(1247) <= not(inputs(123));
    layer0_outputs(1248) <= (inputs(243)) and not (inputs(209));
    layer0_outputs(1249) <= (inputs(162)) and not (inputs(67));
    layer0_outputs(1250) <= not((inputs(192)) or (inputs(151)));
    layer0_outputs(1251) <= not((inputs(41)) xor (inputs(243)));
    layer0_outputs(1252) <= (inputs(40)) or (inputs(55));
    layer0_outputs(1253) <= inputs(119);
    layer0_outputs(1254) <= not((inputs(17)) and (inputs(243)));
    layer0_outputs(1255) <= (inputs(159)) and not (inputs(68));
    layer0_outputs(1256) <= not((inputs(78)) or (inputs(199)));
    layer0_outputs(1257) <= not((inputs(234)) or (inputs(247)));
    layer0_outputs(1258) <= not((inputs(90)) xor (inputs(65)));
    layer0_outputs(1259) <= not((inputs(33)) or (inputs(182)));
    layer0_outputs(1260) <= not((inputs(56)) xor (inputs(252)));
    layer0_outputs(1261) <= not(inputs(100)) or (inputs(23));
    layer0_outputs(1262) <= (inputs(83)) or (inputs(5));
    layer0_outputs(1263) <= not((inputs(120)) xor (inputs(240)));
    layer0_outputs(1264) <= not(inputs(59)) or (inputs(210));
    layer0_outputs(1265) <= (inputs(50)) or (inputs(56));
    layer0_outputs(1266) <= not((inputs(158)) and (inputs(148)));
    layer0_outputs(1267) <= not((inputs(125)) or (inputs(107)));
    layer0_outputs(1268) <= not(inputs(211)) or (inputs(8));
    layer0_outputs(1269) <= inputs(2);
    layer0_outputs(1270) <= not((inputs(239)) xor (inputs(204)));
    layer0_outputs(1271) <= (inputs(215)) and not (inputs(13));
    layer0_outputs(1272) <= not(inputs(133)) or (inputs(254));
    layer0_outputs(1273) <= inputs(91);
    layer0_outputs(1274) <= not(inputs(169));
    layer0_outputs(1275) <= (inputs(143)) or (inputs(51));
    layer0_outputs(1276) <= (inputs(52)) or (inputs(155));
    layer0_outputs(1277) <= inputs(109);
    layer0_outputs(1278) <= (inputs(115)) or (inputs(139));
    layer0_outputs(1279) <= inputs(171);
    layer0_outputs(1280) <= (inputs(195)) xor (inputs(211));
    layer0_outputs(1281) <= not((inputs(225)) xor (inputs(166)));
    layer0_outputs(1282) <= not((inputs(78)) and (inputs(241)));
    layer0_outputs(1283) <= not(inputs(183)) or (inputs(49));
    layer0_outputs(1284) <= not((inputs(65)) or (inputs(178)));
    layer0_outputs(1285) <= (inputs(42)) and (inputs(231));
    layer0_outputs(1286) <= (inputs(122)) and not (inputs(148));
    layer0_outputs(1287) <= not((inputs(253)) and (inputs(3)));
    layer0_outputs(1288) <= not(inputs(0));
    layer0_outputs(1289) <= (inputs(47)) or (inputs(72));
    layer0_outputs(1290) <= (inputs(210)) or (inputs(196));
    layer0_outputs(1291) <= not((inputs(19)) or (inputs(54)));
    layer0_outputs(1292) <= (inputs(42)) and not (inputs(214));
    layer0_outputs(1293) <= not(inputs(52));
    layer0_outputs(1294) <= not(inputs(237));
    layer0_outputs(1295) <= (inputs(52)) or (inputs(10));
    layer0_outputs(1296) <= (inputs(134)) or (inputs(100));
    layer0_outputs(1297) <= (inputs(4)) or (inputs(39));
    layer0_outputs(1298) <= inputs(131);
    layer0_outputs(1299) <= (inputs(129)) xor (inputs(88));
    layer0_outputs(1300) <= inputs(56);
    layer0_outputs(1301) <= (inputs(188)) and not (inputs(28));
    layer0_outputs(1302) <= not((inputs(185)) xor (inputs(142)));
    layer0_outputs(1303) <= not(inputs(66));
    layer0_outputs(1304) <= not((inputs(10)) or (inputs(202)));
    layer0_outputs(1305) <= not(inputs(23));
    layer0_outputs(1306) <= inputs(201);
    layer0_outputs(1307) <= not((inputs(121)) xor (inputs(81)));
    layer0_outputs(1308) <= (inputs(23)) or (inputs(128));
    layer0_outputs(1309) <= (inputs(39)) and not (inputs(233));
    layer0_outputs(1310) <= (inputs(0)) and not (inputs(176));
    layer0_outputs(1311) <= not((inputs(233)) or (inputs(123)));
    layer0_outputs(1312) <= '0';
    layer0_outputs(1313) <= not((inputs(87)) xor (inputs(207)));
    layer0_outputs(1314) <= not((inputs(197)) or (inputs(21)));
    layer0_outputs(1315) <= not((inputs(3)) xor (inputs(234)));
    layer0_outputs(1316) <= not((inputs(165)) or (inputs(234)));
    layer0_outputs(1317) <= inputs(41);
    layer0_outputs(1318) <= not(inputs(118));
    layer0_outputs(1319) <= (inputs(169)) and not (inputs(193));
    layer0_outputs(1320) <= (inputs(120)) or (inputs(166));
    layer0_outputs(1321) <= (inputs(226)) and not (inputs(163));
    layer0_outputs(1322) <= not(inputs(190));
    layer0_outputs(1323) <= not(inputs(216));
    layer0_outputs(1324) <= not(inputs(170));
    layer0_outputs(1325) <= not((inputs(61)) or (inputs(172)));
    layer0_outputs(1326) <= (inputs(224)) and not (inputs(5));
    layer0_outputs(1327) <= not(inputs(105));
    layer0_outputs(1328) <= not((inputs(206)) and (inputs(240)));
    layer0_outputs(1329) <= not((inputs(32)) and (inputs(66)));
    layer0_outputs(1330) <= (inputs(78)) or (inputs(239));
    layer0_outputs(1331) <= (inputs(26)) and not (inputs(241));
    layer0_outputs(1332) <= not((inputs(207)) or (inputs(18)));
    layer0_outputs(1333) <= not(inputs(117));
    layer0_outputs(1334) <= not((inputs(92)) or (inputs(61)));
    layer0_outputs(1335) <= not((inputs(11)) xor (inputs(145)));
    layer0_outputs(1336) <= not(inputs(61));
    layer0_outputs(1337) <= (inputs(166)) and not (inputs(16));
    layer0_outputs(1338) <= inputs(44);
    layer0_outputs(1339) <= (inputs(70)) and not (inputs(34));
    layer0_outputs(1340) <= not(inputs(237));
    layer0_outputs(1341) <= not((inputs(118)) or (inputs(124)));
    layer0_outputs(1342) <= not(inputs(176)) or (inputs(66));
    layer0_outputs(1343) <= (inputs(79)) xor (inputs(185));
    layer0_outputs(1344) <= not((inputs(255)) xor (inputs(217)));
    layer0_outputs(1345) <= inputs(223);
    layer0_outputs(1346) <= not(inputs(117));
    layer0_outputs(1347) <= (inputs(109)) or (inputs(68));
    layer0_outputs(1348) <= not(inputs(72));
    layer0_outputs(1349) <= inputs(160);
    layer0_outputs(1350) <= inputs(60);
    layer0_outputs(1351) <= not(inputs(46));
    layer0_outputs(1352) <= (inputs(175)) xor (inputs(188));
    layer0_outputs(1353) <= (inputs(141)) xor (inputs(113));
    layer0_outputs(1354) <= (inputs(190)) or (inputs(73));
    layer0_outputs(1355) <= not(inputs(217));
    layer0_outputs(1356) <= (inputs(102)) and not (inputs(69));
    layer0_outputs(1357) <= inputs(133);
    layer0_outputs(1358) <= not(inputs(93));
    layer0_outputs(1359) <= not(inputs(137)) or (inputs(45));
    layer0_outputs(1360) <= not((inputs(135)) or (inputs(129)));
    layer0_outputs(1361) <= not(inputs(181));
    layer0_outputs(1362) <= not(inputs(167));
    layer0_outputs(1363) <= not(inputs(130));
    layer0_outputs(1364) <= not((inputs(37)) xor (inputs(238)));
    layer0_outputs(1365) <= (inputs(251)) or (inputs(235));
    layer0_outputs(1366) <= not(inputs(94)) or (inputs(237));
    layer0_outputs(1367) <= '1';
    layer0_outputs(1368) <= '1';
    layer0_outputs(1369) <= not((inputs(243)) or (inputs(195)));
    layer0_outputs(1370) <= (inputs(9)) or (inputs(5));
    layer0_outputs(1371) <= not((inputs(105)) xor (inputs(12)));
    layer0_outputs(1372) <= (inputs(127)) and not (inputs(199));
    layer0_outputs(1373) <= (inputs(185)) and not (inputs(106));
    layer0_outputs(1374) <= inputs(173);
    layer0_outputs(1375) <= (inputs(150)) xor (inputs(0));
    layer0_outputs(1376) <= inputs(138);
    layer0_outputs(1377) <= inputs(136);
    layer0_outputs(1378) <= inputs(198);
    layer0_outputs(1379) <= not((inputs(58)) xor (inputs(91)));
    layer0_outputs(1380) <= '0';
    layer0_outputs(1381) <= not((inputs(164)) xor (inputs(248)));
    layer0_outputs(1382) <= (inputs(198)) xor (inputs(12));
    layer0_outputs(1383) <= (inputs(60)) or (inputs(156));
    layer0_outputs(1384) <= (inputs(213)) or (inputs(198));
    layer0_outputs(1385) <= (inputs(187)) and not (inputs(236));
    layer0_outputs(1386) <= (inputs(172)) or (inputs(167));
    layer0_outputs(1387) <= (inputs(140)) and not (inputs(206));
    layer0_outputs(1388) <= not(inputs(224)) or (inputs(238));
    layer0_outputs(1389) <= not((inputs(162)) or (inputs(109)));
    layer0_outputs(1390) <= not(inputs(96)) or (inputs(240));
    layer0_outputs(1391) <= (inputs(115)) or (inputs(183));
    layer0_outputs(1392) <= not(inputs(52)) or (inputs(114));
    layer0_outputs(1393) <= (inputs(35)) or (inputs(183));
    layer0_outputs(1394) <= (inputs(240)) xor (inputs(228));
    layer0_outputs(1395) <= inputs(117);
    layer0_outputs(1396) <= not((inputs(13)) xor (inputs(60)));
    layer0_outputs(1397) <= (inputs(174)) and not (inputs(245));
    layer0_outputs(1398) <= inputs(211);
    layer0_outputs(1399) <= not((inputs(175)) xor (inputs(131)));
    layer0_outputs(1400) <= not((inputs(44)) or (inputs(97)));
    layer0_outputs(1401) <= inputs(167);
    layer0_outputs(1402) <= not(inputs(206));
    layer0_outputs(1403) <= (inputs(202)) and not (inputs(243));
    layer0_outputs(1404) <= (inputs(171)) and not (inputs(114));
    layer0_outputs(1405) <= inputs(232);
    layer0_outputs(1406) <= (inputs(53)) and not (inputs(77));
    layer0_outputs(1407) <= not((inputs(0)) xor (inputs(14)));
    layer0_outputs(1408) <= not(inputs(41));
    layer0_outputs(1409) <= not((inputs(3)) xor (inputs(134)));
    layer0_outputs(1410) <= inputs(132);
    layer0_outputs(1411) <= (inputs(93)) or (inputs(117));
    layer0_outputs(1412) <= not(inputs(148)) or (inputs(251));
    layer0_outputs(1413) <= (inputs(116)) or (inputs(99));
    layer0_outputs(1414) <= (inputs(152)) and not (inputs(62));
    layer0_outputs(1415) <= inputs(215);
    layer0_outputs(1416) <= (inputs(82)) or (inputs(77));
    layer0_outputs(1417) <= not(inputs(149)) or (inputs(62));
    layer0_outputs(1418) <= not((inputs(17)) or (inputs(70)));
    layer0_outputs(1419) <= not(inputs(103)) or (inputs(24));
    layer0_outputs(1420) <= (inputs(167)) xor (inputs(249));
    layer0_outputs(1421) <= not(inputs(196));
    layer0_outputs(1422) <= not((inputs(227)) or (inputs(88)));
    layer0_outputs(1423) <= inputs(211);
    layer0_outputs(1424) <= '0';
    layer0_outputs(1425) <= (inputs(26)) or (inputs(252));
    layer0_outputs(1426) <= inputs(202);
    layer0_outputs(1427) <= inputs(165);
    layer0_outputs(1428) <= (inputs(164)) or (inputs(59));
    layer0_outputs(1429) <= not((inputs(67)) or (inputs(139)));
    layer0_outputs(1430) <= not((inputs(173)) or (inputs(126)));
    layer0_outputs(1431) <= not(inputs(245)) or (inputs(192));
    layer0_outputs(1432) <= not(inputs(121));
    layer0_outputs(1433) <= not(inputs(213));
    layer0_outputs(1434) <= not(inputs(169)) or (inputs(214));
    layer0_outputs(1435) <= not(inputs(188)) or (inputs(141));
    layer0_outputs(1436) <= not(inputs(120));
    layer0_outputs(1437) <= '0';
    layer0_outputs(1438) <= not((inputs(40)) or (inputs(134)));
    layer0_outputs(1439) <= (inputs(152)) and not (inputs(248));
    layer0_outputs(1440) <= inputs(74);
    layer0_outputs(1441) <= (inputs(105)) and not (inputs(203));
    layer0_outputs(1442) <= not((inputs(69)) or (inputs(76)));
    layer0_outputs(1443) <= not(inputs(148));
    layer0_outputs(1444) <= not(inputs(233));
    layer0_outputs(1445) <= inputs(90);
    layer0_outputs(1446) <= (inputs(28)) or (inputs(142));
    layer0_outputs(1447) <= inputs(255);
    layer0_outputs(1448) <= (inputs(249)) and not (inputs(33));
    layer0_outputs(1449) <= not(inputs(177)) or (inputs(130));
    layer0_outputs(1450) <= inputs(183);
    layer0_outputs(1451) <= not(inputs(140));
    layer0_outputs(1452) <= (inputs(85)) xor (inputs(47));
    layer0_outputs(1453) <= not((inputs(236)) or (inputs(220)));
    layer0_outputs(1454) <= not(inputs(153));
    layer0_outputs(1455) <= (inputs(242)) or (inputs(195));
    layer0_outputs(1456) <= inputs(118);
    layer0_outputs(1457) <= inputs(41);
    layer0_outputs(1458) <= '0';
    layer0_outputs(1459) <= (inputs(85)) or (inputs(96));
    layer0_outputs(1460) <= not(inputs(204));
    layer0_outputs(1461) <= (inputs(115)) and not (inputs(28));
    layer0_outputs(1462) <= (inputs(218)) or (inputs(134));
    layer0_outputs(1463) <= (inputs(238)) xor (inputs(231));
    layer0_outputs(1464) <= not((inputs(11)) or (inputs(231)));
    layer0_outputs(1465) <= not(inputs(238)) or (inputs(29));
    layer0_outputs(1466) <= (inputs(101)) and not (inputs(177));
    layer0_outputs(1467) <= not(inputs(56)) or (inputs(242));
    layer0_outputs(1468) <= (inputs(221)) or (inputs(196));
    layer0_outputs(1469) <= not(inputs(99)) or (inputs(8));
    layer0_outputs(1470) <= (inputs(51)) or (inputs(67));
    layer0_outputs(1471) <= (inputs(90)) and not (inputs(94));
    layer0_outputs(1472) <= not(inputs(215));
    layer0_outputs(1473) <= (inputs(137)) xor (inputs(28));
    layer0_outputs(1474) <= inputs(231);
    layer0_outputs(1475) <= not((inputs(117)) xor (inputs(95)));
    layer0_outputs(1476) <= (inputs(41)) and not (inputs(61));
    layer0_outputs(1477) <= not(inputs(124));
    layer0_outputs(1478) <= (inputs(218)) and not (inputs(198));
    layer0_outputs(1479) <= not(inputs(20)) or (inputs(80));
    layer0_outputs(1480) <= not((inputs(79)) xor (inputs(235)));
    layer0_outputs(1481) <= (inputs(55)) or (inputs(183));
    layer0_outputs(1482) <= (inputs(107)) xor (inputs(190));
    layer0_outputs(1483) <= (inputs(58)) and not (inputs(205));
    layer0_outputs(1484) <= inputs(27);
    layer0_outputs(1485) <= (inputs(218)) and not (inputs(75));
    layer0_outputs(1486) <= '0';
    layer0_outputs(1487) <= (inputs(40)) and not (inputs(117));
    layer0_outputs(1488) <= (inputs(76)) and not (inputs(20));
    layer0_outputs(1489) <= not(inputs(28));
    layer0_outputs(1490) <= not(inputs(6));
    layer0_outputs(1491) <= inputs(163);
    layer0_outputs(1492) <= inputs(224);
    layer0_outputs(1493) <= (inputs(244)) and not (inputs(111));
    layer0_outputs(1494) <= inputs(117);
    layer0_outputs(1495) <= not(inputs(184));
    layer0_outputs(1496) <= (inputs(59)) and not (inputs(20));
    layer0_outputs(1497) <= not(inputs(56)) or (inputs(192));
    layer0_outputs(1498) <= (inputs(102)) and not (inputs(96));
    layer0_outputs(1499) <= not((inputs(43)) xor (inputs(62)));
    layer0_outputs(1500) <= (inputs(107)) or (inputs(19));
    layer0_outputs(1501) <= (inputs(19)) xor (inputs(205));
    layer0_outputs(1502) <= (inputs(63)) and not (inputs(220));
    layer0_outputs(1503) <= (inputs(182)) and not (inputs(93));
    layer0_outputs(1504) <= (inputs(228)) or (inputs(222));
    layer0_outputs(1505) <= (inputs(27)) xor (inputs(169));
    layer0_outputs(1506) <= inputs(233);
    layer0_outputs(1507) <= (inputs(3)) or (inputs(156));
    layer0_outputs(1508) <= (inputs(252)) and not (inputs(254));
    layer0_outputs(1509) <= not((inputs(97)) xor (inputs(33)));
    layer0_outputs(1510) <= not(inputs(77));
    layer0_outputs(1511) <= (inputs(57)) or (inputs(6));
    layer0_outputs(1512) <= inputs(106);
    layer0_outputs(1513) <= inputs(75);
    layer0_outputs(1514) <= (inputs(230)) or (inputs(98));
    layer0_outputs(1515) <= not((inputs(27)) xor (inputs(105)));
    layer0_outputs(1516) <= not((inputs(207)) or (inputs(65)));
    layer0_outputs(1517) <= not(inputs(216)) or (inputs(109));
    layer0_outputs(1518) <= not((inputs(246)) or (inputs(121)));
    layer0_outputs(1519) <= '0';
    layer0_outputs(1520) <= not((inputs(100)) xor (inputs(96)));
    layer0_outputs(1521) <= not(inputs(133));
    layer0_outputs(1522) <= (inputs(89)) and not (inputs(83));
    layer0_outputs(1523) <= not(inputs(224));
    layer0_outputs(1524) <= '0';
    layer0_outputs(1525) <= not(inputs(170)) or (inputs(246));
    layer0_outputs(1526) <= (inputs(233)) or (inputs(210));
    layer0_outputs(1527) <= inputs(94);
    layer0_outputs(1528) <= (inputs(100)) or (inputs(171));
    layer0_outputs(1529) <= (inputs(216)) xor (inputs(30));
    layer0_outputs(1530) <= (inputs(22)) or (inputs(166));
    layer0_outputs(1531) <= not(inputs(202)) or (inputs(32));
    layer0_outputs(1532) <= not(inputs(154)) or (inputs(2));
    layer0_outputs(1533) <= (inputs(109)) or (inputs(143));
    layer0_outputs(1534) <= not((inputs(37)) or (inputs(139)));
    layer0_outputs(1535) <= not(inputs(235)) or (inputs(23));
    layer0_outputs(1536) <= inputs(109);
    layer0_outputs(1537) <= inputs(132);
    layer0_outputs(1538) <= not(inputs(53)) or (inputs(94));
    layer0_outputs(1539) <= inputs(188);
    layer0_outputs(1540) <= not(inputs(139)) or (inputs(237));
    layer0_outputs(1541) <= not((inputs(46)) and (inputs(25)));
    layer0_outputs(1542) <= not(inputs(61)) or (inputs(253));
    layer0_outputs(1543) <= (inputs(44)) and not (inputs(174));
    layer0_outputs(1544) <= not((inputs(236)) and (inputs(238)));
    layer0_outputs(1545) <= (inputs(57)) and not (inputs(12));
    layer0_outputs(1546) <= inputs(182);
    layer0_outputs(1547) <= not(inputs(91)) or (inputs(210));
    layer0_outputs(1548) <= (inputs(16)) xor (inputs(161));
    layer0_outputs(1549) <= (inputs(202)) or (inputs(235));
    layer0_outputs(1550) <= not(inputs(66));
    layer0_outputs(1551) <= inputs(63);
    layer0_outputs(1552) <= not(inputs(205)) or (inputs(96));
    layer0_outputs(1553) <= not(inputs(251));
    layer0_outputs(1554) <= inputs(74);
    layer0_outputs(1555) <= not(inputs(120));
    layer0_outputs(1556) <= inputs(47);
    layer0_outputs(1557) <= not(inputs(140)) or (inputs(130));
    layer0_outputs(1558) <= not(inputs(178));
    layer0_outputs(1559) <= (inputs(43)) xor (inputs(65));
    layer0_outputs(1560) <= (inputs(2)) and not (inputs(212));
    layer0_outputs(1561) <= not(inputs(163));
    layer0_outputs(1562) <= not((inputs(219)) and (inputs(73)));
    layer0_outputs(1563) <= inputs(182);
    layer0_outputs(1564) <= not((inputs(218)) or (inputs(217)));
    layer0_outputs(1565) <= (inputs(126)) and not (inputs(157));
    layer0_outputs(1566) <= not(inputs(179)) or (inputs(125));
    layer0_outputs(1567) <= not((inputs(181)) or (inputs(237)));
    layer0_outputs(1568) <= not(inputs(146));
    layer0_outputs(1569) <= (inputs(26)) xor (inputs(211));
    layer0_outputs(1570) <= inputs(176);
    layer0_outputs(1571) <= '0';
    layer0_outputs(1572) <= (inputs(75)) or (inputs(54));
    layer0_outputs(1573) <= inputs(253);
    layer0_outputs(1574) <= not(inputs(98));
    layer0_outputs(1575) <= not(inputs(119));
    layer0_outputs(1576) <= not((inputs(146)) xor (inputs(211)));
    layer0_outputs(1577) <= not((inputs(117)) or (inputs(215)));
    layer0_outputs(1578) <= not(inputs(71));
    layer0_outputs(1579) <= (inputs(19)) or (inputs(41));
    layer0_outputs(1580) <= inputs(2);
    layer0_outputs(1581) <= (inputs(118)) or (inputs(173));
    layer0_outputs(1582) <= not(inputs(178)) or (inputs(64));
    layer0_outputs(1583) <= inputs(197);
    layer0_outputs(1584) <= not(inputs(179));
    layer0_outputs(1585) <= inputs(34);
    layer0_outputs(1586) <= (inputs(21)) or (inputs(125));
    layer0_outputs(1587) <= not((inputs(239)) or (inputs(239)));
    layer0_outputs(1588) <= inputs(113);
    layer0_outputs(1589) <= not((inputs(17)) xor (inputs(202)));
    layer0_outputs(1590) <= (inputs(67)) or (inputs(131));
    layer0_outputs(1591) <= (inputs(193)) or (inputs(179));
    layer0_outputs(1592) <= not(inputs(69)) or (inputs(160));
    layer0_outputs(1593) <= inputs(151);
    layer0_outputs(1594) <= (inputs(63)) or (inputs(248));
    layer0_outputs(1595) <= (inputs(26)) and not (inputs(143));
    layer0_outputs(1596) <= not((inputs(147)) or (inputs(165)));
    layer0_outputs(1597) <= not((inputs(222)) or (inputs(120)));
    layer0_outputs(1598) <= not((inputs(147)) or (inputs(205)));
    layer0_outputs(1599) <= inputs(111);
    layer0_outputs(1600) <= not(inputs(159));
    layer0_outputs(1601) <= not(inputs(88)) or (inputs(242));
    layer0_outputs(1602) <= inputs(20);
    layer0_outputs(1603) <= (inputs(209)) xor (inputs(100));
    layer0_outputs(1604) <= '0';
    layer0_outputs(1605) <= not(inputs(90));
    layer0_outputs(1606) <= (inputs(0)) and not (inputs(250));
    layer0_outputs(1607) <= not((inputs(158)) xor (inputs(148)));
    layer0_outputs(1608) <= not(inputs(99));
    layer0_outputs(1609) <= not((inputs(174)) xor (inputs(253)));
    layer0_outputs(1610) <= (inputs(201)) and not (inputs(234));
    layer0_outputs(1611) <= not(inputs(99)) or (inputs(153));
    layer0_outputs(1612) <= inputs(117);
    layer0_outputs(1613) <= (inputs(130)) or (inputs(115));
    layer0_outputs(1614) <= '0';
    layer0_outputs(1615) <= '0';
    layer0_outputs(1616) <= not((inputs(141)) or (inputs(140)));
    layer0_outputs(1617) <= inputs(22);
    layer0_outputs(1618) <= not((inputs(241)) xor (inputs(149)));
    layer0_outputs(1619) <= (inputs(57)) and not (inputs(147));
    layer0_outputs(1620) <= not(inputs(182)) or (inputs(60));
    layer0_outputs(1621) <= (inputs(247)) and not (inputs(192));
    layer0_outputs(1622) <= (inputs(133)) or (inputs(175));
    layer0_outputs(1623) <= not(inputs(18));
    layer0_outputs(1624) <= not(inputs(178)) or (inputs(128));
    layer0_outputs(1625) <= inputs(106);
    layer0_outputs(1626) <= not(inputs(213)) or (inputs(41));
    layer0_outputs(1627) <= not(inputs(121));
    layer0_outputs(1628) <= not(inputs(69)) or (inputs(161));
    layer0_outputs(1629) <= (inputs(169)) and not (inputs(252));
    layer0_outputs(1630) <= not((inputs(64)) or (inputs(62)));
    layer0_outputs(1631) <= not(inputs(45));
    layer0_outputs(1632) <= (inputs(126)) or (inputs(152));
    layer0_outputs(1633) <= (inputs(183)) and not (inputs(172));
    layer0_outputs(1634) <= not((inputs(157)) or (inputs(35)));
    layer0_outputs(1635) <= (inputs(135)) and (inputs(198));
    layer0_outputs(1636) <= not((inputs(248)) and (inputs(158)));
    layer0_outputs(1637) <= inputs(38);
    layer0_outputs(1638) <= (inputs(48)) and not (inputs(80));
    layer0_outputs(1639) <= inputs(63);
    layer0_outputs(1640) <= not(inputs(167));
    layer0_outputs(1641) <= not(inputs(127));
    layer0_outputs(1642) <= not((inputs(216)) and (inputs(217)));
    layer0_outputs(1643) <= (inputs(15)) or (inputs(120));
    layer0_outputs(1644) <= not((inputs(22)) xor (inputs(167)));
    layer0_outputs(1645) <= not((inputs(236)) or (inputs(232)));
    layer0_outputs(1646) <= not((inputs(53)) xor (inputs(21)));
    layer0_outputs(1647) <= (inputs(204)) or (inputs(86));
    layer0_outputs(1648) <= (inputs(210)) and not (inputs(64));
    layer0_outputs(1649) <= not((inputs(4)) and (inputs(117)));
    layer0_outputs(1650) <= not(inputs(141));
    layer0_outputs(1651) <= (inputs(136)) and not (inputs(228));
    layer0_outputs(1652) <= not(inputs(75)) or (inputs(221));
    layer0_outputs(1653) <= (inputs(85)) or (inputs(7));
    layer0_outputs(1654) <= inputs(180);
    layer0_outputs(1655) <= not((inputs(94)) or (inputs(109)));
    layer0_outputs(1656) <= '0';
    layer0_outputs(1657) <= not(inputs(108));
    layer0_outputs(1658) <= (inputs(57)) or (inputs(155));
    layer0_outputs(1659) <= not((inputs(209)) or (inputs(127)));
    layer0_outputs(1660) <= not(inputs(43));
    layer0_outputs(1661) <= not(inputs(66)) or (inputs(51));
    layer0_outputs(1662) <= (inputs(233)) and not (inputs(21));
    layer0_outputs(1663) <= not(inputs(104)) or (inputs(99));
    layer0_outputs(1664) <= inputs(108);
    layer0_outputs(1665) <= not((inputs(190)) or (inputs(73)));
    layer0_outputs(1666) <= not((inputs(204)) or (inputs(48)));
    layer0_outputs(1667) <= not((inputs(177)) or (inputs(40)));
    layer0_outputs(1668) <= not(inputs(135));
    layer0_outputs(1669) <= (inputs(75)) or (inputs(55));
    layer0_outputs(1670) <= (inputs(4)) xor (inputs(38));
    layer0_outputs(1671) <= (inputs(188)) xor (inputs(242));
    layer0_outputs(1672) <= (inputs(214)) or (inputs(79));
    layer0_outputs(1673) <= not((inputs(186)) or (inputs(172)));
    layer0_outputs(1674) <= not((inputs(138)) or (inputs(4)));
    layer0_outputs(1675) <= not((inputs(168)) or (inputs(253)));
    layer0_outputs(1676) <= not((inputs(24)) or (inputs(154)));
    layer0_outputs(1677) <= (inputs(113)) or (inputs(83));
    layer0_outputs(1678) <= (inputs(177)) or (inputs(0));
    layer0_outputs(1679) <= (inputs(1)) xor (inputs(145));
    layer0_outputs(1680) <= (inputs(105)) xor (inputs(48));
    layer0_outputs(1681) <= inputs(71);
    layer0_outputs(1682) <= not(inputs(54));
    layer0_outputs(1683) <= inputs(197);
    layer0_outputs(1684) <= not((inputs(162)) or (inputs(32)));
    layer0_outputs(1685) <= (inputs(230)) and not (inputs(211));
    layer0_outputs(1686) <= (inputs(57)) and not (inputs(45));
    layer0_outputs(1687) <= not((inputs(95)) or (inputs(8)));
    layer0_outputs(1688) <= (inputs(232)) and not (inputs(218));
    layer0_outputs(1689) <= not(inputs(197)) or (inputs(10));
    layer0_outputs(1690) <= (inputs(245)) or (inputs(180));
    layer0_outputs(1691) <= (inputs(200)) xor (inputs(248));
    layer0_outputs(1692) <= not(inputs(89));
    layer0_outputs(1693) <= (inputs(29)) xor (inputs(135));
    layer0_outputs(1694) <= (inputs(74)) and not (inputs(194));
    layer0_outputs(1695) <= inputs(86);
    layer0_outputs(1696) <= (inputs(184)) and not (inputs(251));
    layer0_outputs(1697) <= not(inputs(93)) or (inputs(38));
    layer0_outputs(1698) <= (inputs(85)) and not (inputs(188));
    layer0_outputs(1699) <= (inputs(186)) and not (inputs(236));
    layer0_outputs(1700) <= '1';
    layer0_outputs(1701) <= inputs(20);
    layer0_outputs(1702) <= (inputs(21)) or (inputs(27));
    layer0_outputs(1703) <= (inputs(122)) and not (inputs(110));
    layer0_outputs(1704) <= inputs(151);
    layer0_outputs(1705) <= not((inputs(218)) or (inputs(77)));
    layer0_outputs(1706) <= not((inputs(219)) or (inputs(96)));
    layer0_outputs(1707) <= not(inputs(88)) or (inputs(78));
    layer0_outputs(1708) <= (inputs(190)) xor (inputs(15));
    layer0_outputs(1709) <= (inputs(90)) and not (inputs(160));
    layer0_outputs(1710) <= not(inputs(167));
    layer0_outputs(1711) <= (inputs(95)) or (inputs(152));
    layer0_outputs(1712) <= inputs(123);
    layer0_outputs(1713) <= not(inputs(55));
    layer0_outputs(1714) <= not((inputs(16)) and (inputs(190)));
    layer0_outputs(1715) <= (inputs(150)) or (inputs(18));
    layer0_outputs(1716) <= not((inputs(190)) or (inputs(205)));
    layer0_outputs(1717) <= (inputs(1)) xor (inputs(42));
    layer0_outputs(1718) <= not(inputs(217));
    layer0_outputs(1719) <= '1';
    layer0_outputs(1720) <= not(inputs(102)) or (inputs(230));
    layer0_outputs(1721) <= (inputs(195)) and not (inputs(44));
    layer0_outputs(1722) <= inputs(182);
    layer0_outputs(1723) <= not(inputs(99));
    layer0_outputs(1724) <= not((inputs(102)) or (inputs(115)));
    layer0_outputs(1725) <= '0';
    layer0_outputs(1726) <= not((inputs(16)) xor (inputs(0)));
    layer0_outputs(1727) <= (inputs(91)) or (inputs(0));
    layer0_outputs(1728) <= not(inputs(105));
    layer0_outputs(1729) <= (inputs(53)) or (inputs(15));
    layer0_outputs(1730) <= (inputs(44)) or (inputs(113));
    layer0_outputs(1731) <= not((inputs(243)) and (inputs(229)));
    layer0_outputs(1732) <= not(inputs(173));
    layer0_outputs(1733) <= not(inputs(68)) or (inputs(204));
    layer0_outputs(1734) <= inputs(43);
    layer0_outputs(1735) <= not(inputs(221));
    layer0_outputs(1736) <= not(inputs(121)) or (inputs(55));
    layer0_outputs(1737) <= inputs(212);
    layer0_outputs(1738) <= not(inputs(129)) or (inputs(241));
    layer0_outputs(1739) <= inputs(63);
    layer0_outputs(1740) <= not(inputs(49));
    layer0_outputs(1741) <= (inputs(25)) and not (inputs(83));
    layer0_outputs(1742) <= not((inputs(16)) or (inputs(46)));
    layer0_outputs(1743) <= '1';
    layer0_outputs(1744) <= not((inputs(104)) or (inputs(153)));
    layer0_outputs(1745) <= not(inputs(103)) or (inputs(220));
    layer0_outputs(1746) <= (inputs(192)) and not (inputs(47));
    layer0_outputs(1747) <= (inputs(24)) and not (inputs(223));
    layer0_outputs(1748) <= (inputs(245)) and not (inputs(81));
    layer0_outputs(1749) <= not(inputs(116)) or (inputs(244));
    layer0_outputs(1750) <= not((inputs(187)) xor (inputs(66)));
    layer0_outputs(1751) <= not(inputs(165));
    layer0_outputs(1752) <= not(inputs(54)) or (inputs(233));
    layer0_outputs(1753) <= not((inputs(249)) xor (inputs(62)));
    layer0_outputs(1754) <= (inputs(49)) and not (inputs(255));
    layer0_outputs(1755) <= '0';
    layer0_outputs(1756) <= (inputs(5)) and not (inputs(111));
    layer0_outputs(1757) <= inputs(109);
    layer0_outputs(1758) <= (inputs(35)) and not (inputs(250));
    layer0_outputs(1759) <= not((inputs(219)) or (inputs(46)));
    layer0_outputs(1760) <= (inputs(99)) and not (inputs(34));
    layer0_outputs(1761) <= not((inputs(31)) or (inputs(97)));
    layer0_outputs(1762) <= (inputs(105)) or (inputs(80));
    layer0_outputs(1763) <= not((inputs(147)) or (inputs(231)));
    layer0_outputs(1764) <= not((inputs(28)) or (inputs(100)));
    layer0_outputs(1765) <= inputs(41);
    layer0_outputs(1766) <= not((inputs(224)) or (inputs(100)));
    layer0_outputs(1767) <= (inputs(34)) xor (inputs(220));
    layer0_outputs(1768) <= (inputs(33)) or (inputs(197));
    layer0_outputs(1769) <= not(inputs(169));
    layer0_outputs(1770) <= not(inputs(148));
    layer0_outputs(1771) <= not((inputs(165)) or (inputs(0)));
    layer0_outputs(1772) <= not(inputs(160)) or (inputs(228));
    layer0_outputs(1773) <= not(inputs(232)) or (inputs(7));
    layer0_outputs(1774) <= (inputs(84)) and not (inputs(3));
    layer0_outputs(1775) <= not((inputs(181)) or (inputs(157)));
    layer0_outputs(1776) <= inputs(116);
    layer0_outputs(1777) <= not((inputs(76)) xor (inputs(253)));
    layer0_outputs(1778) <= (inputs(58)) or (inputs(51));
    layer0_outputs(1779) <= not(inputs(68)) or (inputs(221));
    layer0_outputs(1780) <= (inputs(201)) and not (inputs(96));
    layer0_outputs(1781) <= not((inputs(168)) or (inputs(69)));
    layer0_outputs(1782) <= (inputs(38)) or (inputs(142));
    layer0_outputs(1783) <= not(inputs(156));
    layer0_outputs(1784) <= '0';
    layer0_outputs(1785) <= not((inputs(240)) and (inputs(209)));
    layer0_outputs(1786) <= (inputs(224)) or (inputs(135));
    layer0_outputs(1787) <= not(inputs(165)) or (inputs(230));
    layer0_outputs(1788) <= not(inputs(190));
    layer0_outputs(1789) <= (inputs(248)) or (inputs(222));
    layer0_outputs(1790) <= not(inputs(238)) or (inputs(254));
    layer0_outputs(1791) <= (inputs(159)) and not (inputs(229));
    layer0_outputs(1792) <= not((inputs(29)) or (inputs(134)));
    layer0_outputs(1793) <= not(inputs(212)) or (inputs(95));
    layer0_outputs(1794) <= '0';
    layer0_outputs(1795) <= (inputs(186)) or (inputs(154));
    layer0_outputs(1796) <= not(inputs(4));
    layer0_outputs(1797) <= not(inputs(57)) or (inputs(234));
    layer0_outputs(1798) <= not(inputs(151)) or (inputs(155));
    layer0_outputs(1799) <= (inputs(46)) or (inputs(8));
    layer0_outputs(1800) <= not(inputs(73));
    layer0_outputs(1801) <= '0';
    layer0_outputs(1802) <= (inputs(36)) xor (inputs(238));
    layer0_outputs(1803) <= inputs(39);
    layer0_outputs(1804) <= (inputs(156)) and not (inputs(34));
    layer0_outputs(1805) <= not((inputs(236)) and (inputs(108)));
    layer0_outputs(1806) <= not(inputs(86));
    layer0_outputs(1807) <= (inputs(209)) or (inputs(195));
    layer0_outputs(1808) <= (inputs(123)) and not (inputs(35));
    layer0_outputs(1809) <= inputs(115);
    layer0_outputs(1810) <= not((inputs(144)) or (inputs(53)));
    layer0_outputs(1811) <= inputs(120);
    layer0_outputs(1812) <= not(inputs(231));
    layer0_outputs(1813) <= not((inputs(58)) or (inputs(180)));
    layer0_outputs(1814) <= '0';
    layer0_outputs(1815) <= (inputs(144)) or (inputs(183));
    layer0_outputs(1816) <= inputs(152);
    layer0_outputs(1817) <= not(inputs(151)) or (inputs(38));
    layer0_outputs(1818) <= (inputs(162)) or (inputs(214));
    layer0_outputs(1819) <= (inputs(55)) or (inputs(209));
    layer0_outputs(1820) <= (inputs(114)) or (inputs(72));
    layer0_outputs(1821) <= not(inputs(106));
    layer0_outputs(1822) <= (inputs(26)) and not (inputs(9));
    layer0_outputs(1823) <= not(inputs(242)) or (inputs(43));
    layer0_outputs(1824) <= (inputs(14)) or (inputs(203));
    layer0_outputs(1825) <= not(inputs(62)) or (inputs(98));
    layer0_outputs(1826) <= not((inputs(222)) xor (inputs(62)));
    layer0_outputs(1827) <= inputs(217);
    layer0_outputs(1828) <= not((inputs(253)) or (inputs(27)));
    layer0_outputs(1829) <= (inputs(192)) and (inputs(79));
    layer0_outputs(1830) <= inputs(152);
    layer0_outputs(1831) <= '0';
    layer0_outputs(1832) <= not(inputs(229)) or (inputs(67));
    layer0_outputs(1833) <= not(inputs(72));
    layer0_outputs(1834) <= not(inputs(56)) or (inputs(216));
    layer0_outputs(1835) <= not(inputs(179)) or (inputs(119));
    layer0_outputs(1836) <= not(inputs(198));
    layer0_outputs(1837) <= inputs(70);
    layer0_outputs(1838) <= (inputs(85)) or (inputs(24));
    layer0_outputs(1839) <= '1';
    layer0_outputs(1840) <= not((inputs(165)) or (inputs(93)));
    layer0_outputs(1841) <= not((inputs(140)) xor (inputs(226)));
    layer0_outputs(1842) <= not((inputs(29)) xor (inputs(125)));
    layer0_outputs(1843) <= (inputs(82)) or (inputs(134));
    layer0_outputs(1844) <= inputs(168);
    layer0_outputs(1845) <= not(inputs(202)) or (inputs(174));
    layer0_outputs(1846) <= (inputs(101)) or (inputs(242));
    layer0_outputs(1847) <= (inputs(181)) and not (inputs(45));
    layer0_outputs(1848) <= not((inputs(212)) xor (inputs(222)));
    layer0_outputs(1849) <= (inputs(66)) and not (inputs(139));
    layer0_outputs(1850) <= not(inputs(52)) or (inputs(124));
    layer0_outputs(1851) <= (inputs(212)) or (inputs(73));
    layer0_outputs(1852) <= inputs(184);
    layer0_outputs(1853) <= (inputs(249)) xor (inputs(226));
    layer0_outputs(1854) <= (inputs(231)) and not (inputs(197));
    layer0_outputs(1855) <= not((inputs(248)) or (inputs(123)));
    layer0_outputs(1856) <= not(inputs(106)) or (inputs(163));
    layer0_outputs(1857) <= (inputs(241)) or (inputs(240));
    layer0_outputs(1858) <= (inputs(185)) xor (inputs(73));
    layer0_outputs(1859) <= not(inputs(85)) or (inputs(218));
    layer0_outputs(1860) <= inputs(22);
    layer0_outputs(1861) <= (inputs(94)) xor (inputs(29));
    layer0_outputs(1862) <= inputs(88);
    layer0_outputs(1863) <= '0';
    layer0_outputs(1864) <= (inputs(51)) and not (inputs(230));
    layer0_outputs(1865) <= not((inputs(191)) xor (inputs(179)));
    layer0_outputs(1866) <= inputs(54);
    layer0_outputs(1867) <= not((inputs(244)) or (inputs(14)));
    layer0_outputs(1868) <= (inputs(210)) and not (inputs(40));
    layer0_outputs(1869) <= '0';
    layer0_outputs(1870) <= not((inputs(136)) or (inputs(168)));
    layer0_outputs(1871) <= not((inputs(235)) xor (inputs(243)));
    layer0_outputs(1872) <= not(inputs(166));
    layer0_outputs(1873) <= not(inputs(203));
    layer0_outputs(1874) <= not((inputs(71)) xor (inputs(56)));
    layer0_outputs(1875) <= '0';
    layer0_outputs(1876) <= not((inputs(27)) or (inputs(116)));
    layer0_outputs(1877) <= '1';
    layer0_outputs(1878) <= not((inputs(36)) xor (inputs(159)));
    layer0_outputs(1879) <= not(inputs(200));
    layer0_outputs(1880) <= (inputs(131)) and not (inputs(35));
    layer0_outputs(1881) <= not(inputs(67));
    layer0_outputs(1882) <= (inputs(20)) and not (inputs(36));
    layer0_outputs(1883) <= (inputs(77)) or (inputs(207));
    layer0_outputs(1884) <= inputs(92);
    layer0_outputs(1885) <= (inputs(26)) xor (inputs(161));
    layer0_outputs(1886) <= (inputs(102)) xor (inputs(5));
    layer0_outputs(1887) <= not((inputs(28)) or (inputs(39)));
    layer0_outputs(1888) <= inputs(119);
    layer0_outputs(1889) <= (inputs(90)) xor (inputs(97));
    layer0_outputs(1890) <= (inputs(189)) or (inputs(248));
    layer0_outputs(1891) <= not(inputs(121)) or (inputs(250));
    layer0_outputs(1892) <= not(inputs(52)) or (inputs(16));
    layer0_outputs(1893) <= not((inputs(217)) or (inputs(254)));
    layer0_outputs(1894) <= (inputs(240)) xor (inputs(173));
    layer0_outputs(1895) <= not((inputs(154)) or (inputs(27)));
    layer0_outputs(1896) <= (inputs(137)) and not (inputs(194));
    layer0_outputs(1897) <= inputs(34);
    layer0_outputs(1898) <= (inputs(10)) and not (inputs(128));
    layer0_outputs(1899) <= (inputs(15)) or (inputs(55));
    layer0_outputs(1900) <= not((inputs(71)) or (inputs(1)));
    layer0_outputs(1901) <= not(inputs(53)) or (inputs(10));
    layer0_outputs(1902) <= not(inputs(180)) or (inputs(247));
    layer0_outputs(1903) <= not(inputs(188));
    layer0_outputs(1904) <= not((inputs(135)) xor (inputs(161)));
    layer0_outputs(1905) <= not((inputs(37)) or (inputs(22)));
    layer0_outputs(1906) <= not((inputs(40)) or (inputs(246)));
    layer0_outputs(1907) <= not(inputs(54));
    layer0_outputs(1908) <= not((inputs(23)) or (inputs(124)));
    layer0_outputs(1909) <= (inputs(84)) and not (inputs(173));
    layer0_outputs(1910) <= not((inputs(10)) or (inputs(15)));
    layer0_outputs(1911) <= not(inputs(108)) or (inputs(98));
    layer0_outputs(1912) <= (inputs(216)) and not (inputs(6));
    layer0_outputs(1913) <= inputs(102);
    layer0_outputs(1914) <= (inputs(138)) or (inputs(145));
    layer0_outputs(1915) <= not((inputs(215)) xor (inputs(50)));
    layer0_outputs(1916) <= (inputs(158)) xor (inputs(125));
    layer0_outputs(1917) <= (inputs(178)) or (inputs(21));
    layer0_outputs(1918) <= inputs(197);
    layer0_outputs(1919) <= '0';
    layer0_outputs(1920) <= (inputs(128)) xor (inputs(13));
    layer0_outputs(1921) <= (inputs(245)) or (inputs(100));
    layer0_outputs(1922) <= not((inputs(109)) or (inputs(241)));
    layer0_outputs(1923) <= inputs(24);
    layer0_outputs(1924) <= not((inputs(249)) xor (inputs(196)));
    layer0_outputs(1925) <= not(inputs(151));
    layer0_outputs(1926) <= (inputs(51)) or (inputs(119));
    layer0_outputs(1927) <= (inputs(31)) or (inputs(204));
    layer0_outputs(1928) <= inputs(54);
    layer0_outputs(1929) <= (inputs(41)) xor (inputs(1));
    layer0_outputs(1930) <= not((inputs(79)) and (inputs(98)));
    layer0_outputs(1931) <= (inputs(118)) or (inputs(157));
    layer0_outputs(1932) <= (inputs(200)) or (inputs(174));
    layer0_outputs(1933) <= inputs(167);
    layer0_outputs(1934) <= (inputs(15)) xor (inputs(229));
    layer0_outputs(1935) <= inputs(225);
    layer0_outputs(1936) <= '1';
    layer0_outputs(1937) <= not(inputs(173)) or (inputs(45));
    layer0_outputs(1938) <= not(inputs(55));
    layer0_outputs(1939) <= not(inputs(175)) or (inputs(64));
    layer0_outputs(1940) <= (inputs(162)) and not (inputs(238));
    layer0_outputs(1941) <= (inputs(144)) or (inputs(61));
    layer0_outputs(1942) <= not((inputs(46)) xor (inputs(235)));
    layer0_outputs(1943) <= not((inputs(212)) or (inputs(76)));
    layer0_outputs(1944) <= inputs(141);
    layer0_outputs(1945) <= (inputs(76)) and not (inputs(40));
    layer0_outputs(1946) <= not((inputs(188)) or (inputs(201)));
    layer0_outputs(1947) <= not(inputs(139));
    layer0_outputs(1948) <= not(inputs(183));
    layer0_outputs(1949) <= (inputs(82)) or (inputs(85));
    layer0_outputs(1950) <= inputs(189);
    layer0_outputs(1951) <= not(inputs(124));
    layer0_outputs(1952) <= (inputs(34)) and (inputs(184));
    layer0_outputs(1953) <= (inputs(58)) xor (inputs(66));
    layer0_outputs(1954) <= (inputs(167)) and not (inputs(115));
    layer0_outputs(1955) <= not((inputs(245)) xor (inputs(25)));
    layer0_outputs(1956) <= inputs(164);
    layer0_outputs(1957) <= (inputs(26)) xor (inputs(150));
    layer0_outputs(1958) <= not(inputs(20)) or (inputs(43));
    layer0_outputs(1959) <= inputs(164);
    layer0_outputs(1960) <= (inputs(37)) xor (inputs(77));
    layer0_outputs(1961) <= (inputs(150)) or (inputs(127));
    layer0_outputs(1962) <= not(inputs(87)) or (inputs(3));
    layer0_outputs(1963) <= not(inputs(101));
    layer0_outputs(1964) <= (inputs(157)) or (inputs(228));
    layer0_outputs(1965) <= not((inputs(23)) xor (inputs(207)));
    layer0_outputs(1966) <= inputs(201);
    layer0_outputs(1967) <= not(inputs(125)) or (inputs(234));
    layer0_outputs(1968) <= not((inputs(83)) or (inputs(53)));
    layer0_outputs(1969) <= (inputs(138)) or (inputs(172));
    layer0_outputs(1970) <= (inputs(245)) or (inputs(157));
    layer0_outputs(1971) <= (inputs(206)) or (inputs(196));
    layer0_outputs(1972) <= not(inputs(62));
    layer0_outputs(1973) <= not(inputs(213));
    layer0_outputs(1974) <= not(inputs(179));
    layer0_outputs(1975) <= not((inputs(137)) xor (inputs(114)));
    layer0_outputs(1976) <= (inputs(95)) xor (inputs(222));
    layer0_outputs(1977) <= inputs(218);
    layer0_outputs(1978) <= (inputs(101)) xor (inputs(87));
    layer0_outputs(1979) <= inputs(216);
    layer0_outputs(1980) <= not((inputs(84)) or (inputs(246)));
    layer0_outputs(1981) <= not(inputs(112));
    layer0_outputs(1982) <= inputs(199);
    layer0_outputs(1983) <= not((inputs(31)) xor (inputs(229)));
    layer0_outputs(1984) <= (inputs(132)) and not (inputs(179));
    layer0_outputs(1985) <= not(inputs(184)) or (inputs(232));
    layer0_outputs(1986) <= not(inputs(172)) or (inputs(16));
    layer0_outputs(1987) <= not((inputs(62)) or (inputs(147)));
    layer0_outputs(1988) <= (inputs(50)) and (inputs(37));
    layer0_outputs(1989) <= inputs(52);
    layer0_outputs(1990) <= not(inputs(113)) or (inputs(130));
    layer0_outputs(1991) <= not((inputs(185)) xor (inputs(5)));
    layer0_outputs(1992) <= not((inputs(182)) or (inputs(111)));
    layer0_outputs(1993) <= (inputs(166)) or (inputs(168));
    layer0_outputs(1994) <= not((inputs(164)) or (inputs(221)));
    layer0_outputs(1995) <= '0';
    layer0_outputs(1996) <= not(inputs(148));
    layer0_outputs(1997) <= not(inputs(149));
    layer0_outputs(1998) <= not(inputs(141)) or (inputs(47));
    layer0_outputs(1999) <= (inputs(13)) xor (inputs(107));
    layer0_outputs(2000) <= (inputs(84)) xor (inputs(252));
    layer0_outputs(2001) <= inputs(143);
    layer0_outputs(2002) <= not(inputs(252));
    layer0_outputs(2003) <= not((inputs(95)) xor (inputs(197)));
    layer0_outputs(2004) <= (inputs(36)) or (inputs(174));
    layer0_outputs(2005) <= (inputs(122)) and not (inputs(213));
    layer0_outputs(2006) <= inputs(152);
    layer0_outputs(2007) <= not((inputs(107)) or (inputs(31)));
    layer0_outputs(2008) <= inputs(235);
    layer0_outputs(2009) <= not(inputs(172));
    layer0_outputs(2010) <= inputs(214);
    layer0_outputs(2011) <= not((inputs(198)) or (inputs(92)));
    layer0_outputs(2012) <= not((inputs(39)) or (inputs(22)));
    layer0_outputs(2013) <= inputs(194);
    layer0_outputs(2014) <= (inputs(156)) and not (inputs(98));
    layer0_outputs(2015) <= not((inputs(183)) and (inputs(186)));
    layer0_outputs(2016) <= (inputs(2)) xor (inputs(50));
    layer0_outputs(2017) <= (inputs(208)) and not (inputs(104));
    layer0_outputs(2018) <= not((inputs(214)) or (inputs(61)));
    layer0_outputs(2019) <= inputs(62);
    layer0_outputs(2020) <= (inputs(170)) or (inputs(253));
    layer0_outputs(2021) <= not(inputs(73));
    layer0_outputs(2022) <= inputs(107);
    layer0_outputs(2023) <= not(inputs(156)) or (inputs(225));
    layer0_outputs(2024) <= (inputs(213)) and not (inputs(78));
    layer0_outputs(2025) <= (inputs(87)) and not (inputs(51));
    layer0_outputs(2026) <= not(inputs(232));
    layer0_outputs(2027) <= not((inputs(158)) or (inputs(240)));
    layer0_outputs(2028) <= not((inputs(179)) or (inputs(6)));
    layer0_outputs(2029) <= inputs(181);
    layer0_outputs(2030) <= not(inputs(69)) or (inputs(177));
    layer0_outputs(2031) <= not(inputs(169));
    layer0_outputs(2032) <= not((inputs(62)) xor (inputs(23)));
    layer0_outputs(2033) <= not((inputs(3)) and (inputs(203)));
    layer0_outputs(2034) <= not(inputs(88));
    layer0_outputs(2035) <= not((inputs(99)) and (inputs(223)));
    layer0_outputs(2036) <= inputs(198);
    layer0_outputs(2037) <= not(inputs(118));
    layer0_outputs(2038) <= not(inputs(144)) or (inputs(160));
    layer0_outputs(2039) <= (inputs(230)) and not (inputs(196));
    layer0_outputs(2040) <= not(inputs(156));
    layer0_outputs(2041) <= inputs(132);
    layer0_outputs(2042) <= not((inputs(114)) or (inputs(133)));
    layer0_outputs(2043) <= (inputs(217)) and not (inputs(108));
    layer0_outputs(2044) <= not(inputs(137));
    layer0_outputs(2045) <= not((inputs(78)) or (inputs(165)));
    layer0_outputs(2046) <= (inputs(36)) or (inputs(27));
    layer0_outputs(2047) <= not((inputs(7)) xor (inputs(52)));
    layer0_outputs(2048) <= not(inputs(127));
    layer0_outputs(2049) <= not((inputs(122)) or (inputs(160)));
    layer0_outputs(2050) <= (inputs(224)) xor (inputs(11));
    layer0_outputs(2051) <= not((inputs(34)) and (inputs(111)));
    layer0_outputs(2052) <= inputs(181);
    layer0_outputs(2053) <= (inputs(20)) and not (inputs(130));
    layer0_outputs(2054) <= (inputs(164)) and not (inputs(98));
    layer0_outputs(2055) <= not((inputs(54)) or (inputs(120)));
    layer0_outputs(2056) <= (inputs(158)) or (inputs(245));
    layer0_outputs(2057) <= (inputs(123)) and not (inputs(7));
    layer0_outputs(2058) <= inputs(218);
    layer0_outputs(2059) <= not((inputs(170)) xor (inputs(76)));
    layer0_outputs(2060) <= (inputs(167)) and not (inputs(5));
    layer0_outputs(2061) <= (inputs(64)) and not (inputs(32));
    layer0_outputs(2062) <= (inputs(97)) and not (inputs(16));
    layer0_outputs(2063) <= (inputs(171)) and not (inputs(240));
    layer0_outputs(2064) <= not(inputs(210));
    layer0_outputs(2065) <= inputs(185);
    layer0_outputs(2066) <= not((inputs(237)) or (inputs(239)));
    layer0_outputs(2067) <= inputs(75);
    layer0_outputs(2068) <= (inputs(127)) xor (inputs(103));
    layer0_outputs(2069) <= (inputs(228)) or (inputs(129));
    layer0_outputs(2070) <= inputs(83);
    layer0_outputs(2071) <= not(inputs(165)) or (inputs(216));
    layer0_outputs(2072) <= (inputs(8)) xor (inputs(254));
    layer0_outputs(2073) <= inputs(151);
    layer0_outputs(2074) <= (inputs(194)) and not (inputs(207));
    layer0_outputs(2075) <= not((inputs(95)) xor (inputs(134)));
    layer0_outputs(2076) <= inputs(161);
    layer0_outputs(2077) <= not((inputs(211)) or (inputs(244)));
    layer0_outputs(2078) <= not((inputs(30)) and (inputs(223)));
    layer0_outputs(2079) <= not(inputs(241));
    layer0_outputs(2080) <= not((inputs(99)) or (inputs(61)));
    layer0_outputs(2081) <= not((inputs(241)) and (inputs(4)));
    layer0_outputs(2082) <= (inputs(2)) and not (inputs(17));
    layer0_outputs(2083) <= not((inputs(12)) xor (inputs(76)));
    layer0_outputs(2084) <= not(inputs(75));
    layer0_outputs(2085) <= not((inputs(253)) or (inputs(154)));
    layer0_outputs(2086) <= not((inputs(109)) xor (inputs(254)));
    layer0_outputs(2087) <= (inputs(186)) or (inputs(70));
    layer0_outputs(2088) <= (inputs(42)) or (inputs(187));
    layer0_outputs(2089) <= not((inputs(182)) or (inputs(158)));
    layer0_outputs(2090) <= (inputs(13)) or (inputs(209));
    layer0_outputs(2091) <= not(inputs(248)) or (inputs(208));
    layer0_outputs(2092) <= '0';
    layer0_outputs(2093) <= not((inputs(32)) or (inputs(204)));
    layer0_outputs(2094) <= (inputs(38)) and not (inputs(221));
    layer0_outputs(2095) <= inputs(244);
    layer0_outputs(2096) <= inputs(235);
    layer0_outputs(2097) <= not((inputs(83)) xor (inputs(233)));
    layer0_outputs(2098) <= not((inputs(177)) or (inputs(16)));
    layer0_outputs(2099) <= not(inputs(71)) or (inputs(6));
    layer0_outputs(2100) <= not((inputs(214)) or (inputs(19)));
    layer0_outputs(2101) <= (inputs(91)) or (inputs(196));
    layer0_outputs(2102) <= not((inputs(196)) xor (inputs(47)));
    layer0_outputs(2103) <= not((inputs(245)) or (inputs(199)));
    layer0_outputs(2104) <= not(inputs(163));
    layer0_outputs(2105) <= not(inputs(131));
    layer0_outputs(2106) <= (inputs(103)) and not (inputs(234));
    layer0_outputs(2107) <= not((inputs(173)) or (inputs(164)));
    layer0_outputs(2108) <= inputs(108);
    layer0_outputs(2109) <= not(inputs(133)) or (inputs(111));
    layer0_outputs(2110) <= (inputs(151)) and not (inputs(206));
    layer0_outputs(2111) <= (inputs(14)) xor (inputs(45));
    layer0_outputs(2112) <= not(inputs(55)) or (inputs(144));
    layer0_outputs(2113) <= not(inputs(86));
    layer0_outputs(2114) <= inputs(217);
    layer0_outputs(2115) <= not((inputs(115)) or (inputs(44)));
    layer0_outputs(2116) <= not(inputs(162)) or (inputs(98));
    layer0_outputs(2117) <= (inputs(235)) and not (inputs(236));
    layer0_outputs(2118) <= (inputs(156)) and not (inputs(164));
    layer0_outputs(2119) <= (inputs(222)) or (inputs(78));
    layer0_outputs(2120) <= not((inputs(184)) xor (inputs(96)));
    layer0_outputs(2121) <= (inputs(227)) xor (inputs(40));
    layer0_outputs(2122) <= (inputs(42)) or (inputs(68));
    layer0_outputs(2123) <= (inputs(246)) and not (inputs(28));
    layer0_outputs(2124) <= inputs(44);
    layer0_outputs(2125) <= not((inputs(31)) or (inputs(97)));
    layer0_outputs(2126) <= inputs(195);
    layer0_outputs(2127) <= '0';
    layer0_outputs(2128) <= (inputs(145)) xor (inputs(217));
    layer0_outputs(2129) <= (inputs(154)) and not (inputs(79));
    layer0_outputs(2130) <= not((inputs(76)) xor (inputs(51)));
    layer0_outputs(2131) <= not(inputs(71)) or (inputs(11));
    layer0_outputs(2132) <= not((inputs(227)) xor (inputs(100)));
    layer0_outputs(2133) <= not((inputs(103)) or (inputs(103)));
    layer0_outputs(2134) <= not((inputs(201)) or (inputs(155)));
    layer0_outputs(2135) <= (inputs(240)) and (inputs(212));
    layer0_outputs(2136) <= not(inputs(162));
    layer0_outputs(2137) <= (inputs(78)) or (inputs(136));
    layer0_outputs(2138) <= not((inputs(48)) or (inputs(74)));
    layer0_outputs(2139) <= inputs(107);
    layer0_outputs(2140) <= (inputs(246)) and not (inputs(160));
    layer0_outputs(2141) <= not(inputs(146));
    layer0_outputs(2142) <= not(inputs(88));
    layer0_outputs(2143) <= not(inputs(153)) or (inputs(54));
    layer0_outputs(2144) <= not(inputs(76));
    layer0_outputs(2145) <= not(inputs(158));
    layer0_outputs(2146) <= not(inputs(185)) or (inputs(89));
    layer0_outputs(2147) <= not(inputs(38));
    layer0_outputs(2148) <= not(inputs(103));
    layer0_outputs(2149) <= not(inputs(163));
    layer0_outputs(2150) <= not(inputs(213));
    layer0_outputs(2151) <= not(inputs(46));
    layer0_outputs(2152) <= (inputs(157)) xor (inputs(4));
    layer0_outputs(2153) <= (inputs(17)) xor (inputs(245));
    layer0_outputs(2154) <= (inputs(215)) and not (inputs(21));
    layer0_outputs(2155) <= (inputs(251)) and not (inputs(249));
    layer0_outputs(2156) <= not(inputs(39)) or (inputs(101));
    layer0_outputs(2157) <= inputs(144);
    layer0_outputs(2158) <= '0';
    layer0_outputs(2159) <= inputs(138);
    layer0_outputs(2160) <= not((inputs(227)) or (inputs(210)));
    layer0_outputs(2161) <= not(inputs(237));
    layer0_outputs(2162) <= not(inputs(170)) or (inputs(219));
    layer0_outputs(2163) <= not(inputs(91));
    layer0_outputs(2164) <= not((inputs(8)) and (inputs(247)));
    layer0_outputs(2165) <= '0';
    layer0_outputs(2166) <= (inputs(194)) and not (inputs(243));
    layer0_outputs(2167) <= not(inputs(101));
    layer0_outputs(2168) <= inputs(9);
    layer0_outputs(2169) <= not((inputs(198)) or (inputs(45)));
    layer0_outputs(2170) <= inputs(101);
    layer0_outputs(2171) <= not(inputs(213)) or (inputs(98));
    layer0_outputs(2172) <= not(inputs(116));
    layer0_outputs(2173) <= not(inputs(57));
    layer0_outputs(2174) <= '1';
    layer0_outputs(2175) <= inputs(155);
    layer0_outputs(2176) <= not((inputs(146)) or (inputs(201)));
    layer0_outputs(2177) <= not((inputs(47)) or (inputs(110)));
    layer0_outputs(2178) <= (inputs(83)) xor (inputs(241));
    layer0_outputs(2179) <= (inputs(243)) xor (inputs(75));
    layer0_outputs(2180) <= not((inputs(106)) xor (inputs(49)));
    layer0_outputs(2181) <= '1';
    layer0_outputs(2182) <= not((inputs(86)) or (inputs(125)));
    layer0_outputs(2183) <= not((inputs(9)) or (inputs(16)));
    layer0_outputs(2184) <= '0';
    layer0_outputs(2185) <= (inputs(146)) and not (inputs(46));
    layer0_outputs(2186) <= inputs(153);
    layer0_outputs(2187) <= not(inputs(134));
    layer0_outputs(2188) <= not(inputs(147)) or (inputs(24));
    layer0_outputs(2189) <= not(inputs(36));
    layer0_outputs(2190) <= (inputs(71)) or (inputs(250));
    layer0_outputs(2191) <= (inputs(69)) xor (inputs(140));
    layer0_outputs(2192) <= not((inputs(34)) xor (inputs(156)));
    layer0_outputs(2193) <= (inputs(34)) and (inputs(127));
    layer0_outputs(2194) <= '0';
    layer0_outputs(2195) <= not(inputs(123));
    layer0_outputs(2196) <= not((inputs(179)) or (inputs(187)));
    layer0_outputs(2197) <= (inputs(162)) xor (inputs(3));
    layer0_outputs(2198) <= not(inputs(98));
    layer0_outputs(2199) <= inputs(167);
    layer0_outputs(2200) <= (inputs(190)) or (inputs(202));
    layer0_outputs(2201) <= inputs(255);
    layer0_outputs(2202) <= not(inputs(52));
    layer0_outputs(2203) <= not(inputs(88)) or (inputs(149));
    layer0_outputs(2204) <= (inputs(85)) and (inputs(176));
    layer0_outputs(2205) <= not(inputs(197)) or (inputs(34));
    layer0_outputs(2206) <= (inputs(216)) or (inputs(75));
    layer0_outputs(2207) <= (inputs(31)) xor (inputs(203));
    layer0_outputs(2208) <= not((inputs(238)) and (inputs(147)));
    layer0_outputs(2209) <= not(inputs(220)) or (inputs(30));
    layer0_outputs(2210) <= '1';
    layer0_outputs(2211) <= (inputs(223)) and not (inputs(244));
    layer0_outputs(2212) <= not(inputs(100));
    layer0_outputs(2213) <= not(inputs(220)) or (inputs(245));
    layer0_outputs(2214) <= not((inputs(71)) or (inputs(255)));
    layer0_outputs(2215) <= inputs(93);
    layer0_outputs(2216) <= not((inputs(88)) xor (inputs(160)));
    layer0_outputs(2217) <= not((inputs(41)) or (inputs(130)));
    layer0_outputs(2218) <= '0';
    layer0_outputs(2219) <= not((inputs(184)) or (inputs(28)));
    layer0_outputs(2220) <= (inputs(194)) xor (inputs(94));
    layer0_outputs(2221) <= (inputs(172)) or (inputs(34));
    layer0_outputs(2222) <= inputs(29);
    layer0_outputs(2223) <= not(inputs(39)) or (inputs(250));
    layer0_outputs(2224) <= not((inputs(220)) and (inputs(131)));
    layer0_outputs(2225) <= not(inputs(153)) or (inputs(59));
    layer0_outputs(2226) <= inputs(54);
    layer0_outputs(2227) <= not(inputs(101));
    layer0_outputs(2228) <= not(inputs(65)) or (inputs(83));
    layer0_outputs(2229) <= (inputs(29)) xor (inputs(162));
    layer0_outputs(2230) <= (inputs(126)) xor (inputs(42));
    layer0_outputs(2231) <= not((inputs(169)) xor (inputs(137)));
    layer0_outputs(2232) <= not(inputs(19));
    layer0_outputs(2233) <= (inputs(223)) and not (inputs(181));
    layer0_outputs(2234) <= inputs(138);
    layer0_outputs(2235) <= '1';
    layer0_outputs(2236) <= not((inputs(1)) xor (inputs(75)));
    layer0_outputs(2237) <= not((inputs(144)) and (inputs(249)));
    layer0_outputs(2238) <= (inputs(129)) and not (inputs(108));
    layer0_outputs(2239) <= not((inputs(154)) or (inputs(65)));
    layer0_outputs(2240) <= (inputs(128)) and not (inputs(241));
    layer0_outputs(2241) <= (inputs(226)) or (inputs(35));
    layer0_outputs(2242) <= not((inputs(59)) or (inputs(103)));
    layer0_outputs(2243) <= (inputs(99)) xor (inputs(120));
    layer0_outputs(2244) <= (inputs(172)) or (inputs(204));
    layer0_outputs(2245) <= (inputs(184)) and not (inputs(107));
    layer0_outputs(2246) <= inputs(76);
    layer0_outputs(2247) <= (inputs(216)) and not (inputs(5));
    layer0_outputs(2248) <= not(inputs(90)) or (inputs(89));
    layer0_outputs(2249) <= (inputs(211)) or (inputs(196));
    layer0_outputs(2250) <= not(inputs(72));
    layer0_outputs(2251) <= (inputs(208)) and (inputs(158));
    layer0_outputs(2252) <= (inputs(25)) or (inputs(156));
    layer0_outputs(2253) <= not(inputs(202)) or (inputs(0));
    layer0_outputs(2254) <= not((inputs(12)) xor (inputs(192)));
    layer0_outputs(2255) <= inputs(122);
    layer0_outputs(2256) <= not((inputs(20)) or (inputs(171)));
    layer0_outputs(2257) <= not(inputs(116));
    layer0_outputs(2258) <= not(inputs(148)) or (inputs(29));
    layer0_outputs(2259) <= not((inputs(82)) or (inputs(160)));
    layer0_outputs(2260) <= (inputs(143)) and not (inputs(79));
    layer0_outputs(2261) <= (inputs(215)) and not (inputs(225));
    layer0_outputs(2262) <= (inputs(64)) and not (inputs(175));
    layer0_outputs(2263) <= (inputs(73)) xor (inputs(239));
    layer0_outputs(2264) <= (inputs(99)) or (inputs(175));
    layer0_outputs(2265) <= not((inputs(163)) or (inputs(164)));
    layer0_outputs(2266) <= inputs(148);
    layer0_outputs(2267) <= (inputs(210)) or (inputs(219));
    layer0_outputs(2268) <= (inputs(108)) and not (inputs(112));
    layer0_outputs(2269) <= not((inputs(68)) or (inputs(212)));
    layer0_outputs(2270) <= not(inputs(197));
    layer0_outputs(2271) <= not(inputs(246)) or (inputs(131));
    layer0_outputs(2272) <= (inputs(6)) or (inputs(21));
    layer0_outputs(2273) <= inputs(97);
    layer0_outputs(2274) <= not(inputs(1));
    layer0_outputs(2275) <= not((inputs(179)) xor (inputs(209)));
    layer0_outputs(2276) <= inputs(132);
    layer0_outputs(2277) <= (inputs(77)) and not (inputs(237));
    layer0_outputs(2278) <= inputs(119);
    layer0_outputs(2279) <= not(inputs(37));
    layer0_outputs(2280) <= (inputs(68)) and not (inputs(48));
    layer0_outputs(2281) <= (inputs(142)) xor (inputs(93));
    layer0_outputs(2282) <= (inputs(43)) and not (inputs(253));
    layer0_outputs(2283) <= not((inputs(225)) or (inputs(168)));
    layer0_outputs(2284) <= inputs(165);
    layer0_outputs(2285) <= not((inputs(180)) xor (inputs(205)));
    layer0_outputs(2286) <= not(inputs(112)) or (inputs(84));
    layer0_outputs(2287) <= not(inputs(72)) or (inputs(61));
    layer0_outputs(2288) <= not((inputs(136)) or (inputs(178)));
    layer0_outputs(2289) <= (inputs(206)) or (inputs(188));
    layer0_outputs(2290) <= (inputs(214)) and not (inputs(4));
    layer0_outputs(2291) <= (inputs(123)) or (inputs(230));
    layer0_outputs(2292) <= not(inputs(142));
    layer0_outputs(2293) <= (inputs(67)) and not (inputs(239));
    layer0_outputs(2294) <= not((inputs(154)) or (inputs(134)));
    layer0_outputs(2295) <= not(inputs(151)) or (inputs(80));
    layer0_outputs(2296) <= not((inputs(198)) or (inputs(194)));
    layer0_outputs(2297) <= not(inputs(142));
    layer0_outputs(2298) <= not(inputs(72));
    layer0_outputs(2299) <= not((inputs(162)) or (inputs(145)));
    layer0_outputs(2300) <= not(inputs(56)) or (inputs(27));
    layer0_outputs(2301) <= (inputs(190)) xor (inputs(17));
    layer0_outputs(2302) <= not((inputs(64)) or (inputs(140)));
    layer0_outputs(2303) <= not((inputs(7)) and (inputs(146)));
    layer0_outputs(2304) <= (inputs(231)) and not (inputs(127));
    layer0_outputs(2305) <= not((inputs(110)) xor (inputs(253)));
    layer0_outputs(2306) <= inputs(224);
    layer0_outputs(2307) <= (inputs(182)) xor (inputs(254));
    layer0_outputs(2308) <= (inputs(213)) or (inputs(74));
    layer0_outputs(2309) <= (inputs(51)) or (inputs(49));
    layer0_outputs(2310) <= not((inputs(228)) xor (inputs(113)));
    layer0_outputs(2311) <= not(inputs(119)) or (inputs(12));
    layer0_outputs(2312) <= (inputs(209)) or (inputs(151));
    layer0_outputs(2313) <= '1';
    layer0_outputs(2314) <= not((inputs(133)) and (inputs(133)));
    layer0_outputs(2315) <= inputs(106);
    layer0_outputs(2316) <= (inputs(42)) or (inputs(57));
    layer0_outputs(2317) <= not(inputs(255)) or (inputs(99));
    layer0_outputs(2318) <= (inputs(229)) and not (inputs(175));
    layer0_outputs(2319) <= not(inputs(112)) or (inputs(146));
    layer0_outputs(2320) <= not((inputs(59)) and (inputs(222)));
    layer0_outputs(2321) <= not(inputs(45)) or (inputs(144));
    layer0_outputs(2322) <= not(inputs(152));
    layer0_outputs(2323) <= not(inputs(100)) or (inputs(174));
    layer0_outputs(2324) <= (inputs(191)) and (inputs(184));
    layer0_outputs(2325) <= (inputs(183)) and not (inputs(131));
    layer0_outputs(2326) <= (inputs(21)) or (inputs(186));
    layer0_outputs(2327) <= not((inputs(58)) or (inputs(105)));
    layer0_outputs(2328) <= inputs(236);
    layer0_outputs(2329) <= '0';
    layer0_outputs(2330) <= '0';
    layer0_outputs(2331) <= not(inputs(53)) or (inputs(243));
    layer0_outputs(2332) <= not((inputs(110)) and (inputs(177)));
    layer0_outputs(2333) <= '0';
    layer0_outputs(2334) <= not(inputs(155)) or (inputs(244));
    layer0_outputs(2335) <= (inputs(210)) and not (inputs(251));
    layer0_outputs(2336) <= not((inputs(81)) xor (inputs(151)));
    layer0_outputs(2337) <= (inputs(253)) xor (inputs(50));
    layer0_outputs(2338) <= inputs(61);
    layer0_outputs(2339) <= (inputs(169)) or (inputs(22));
    layer0_outputs(2340) <= '0';
    layer0_outputs(2341) <= (inputs(104)) and (inputs(46));
    layer0_outputs(2342) <= not(inputs(155)) or (inputs(16));
    layer0_outputs(2343) <= not(inputs(96));
    layer0_outputs(2344) <= not(inputs(5)) or (inputs(96));
    layer0_outputs(2345) <= (inputs(242)) or (inputs(100));
    layer0_outputs(2346) <= inputs(132);
    layer0_outputs(2347) <= '0';
    layer0_outputs(2348) <= inputs(150);
    layer0_outputs(2349) <= not(inputs(207));
    layer0_outputs(2350) <= (inputs(195)) or (inputs(198));
    layer0_outputs(2351) <= not((inputs(144)) xor (inputs(224)));
    layer0_outputs(2352) <= not(inputs(199)) or (inputs(130));
    layer0_outputs(2353) <= not(inputs(189));
    layer0_outputs(2354) <= '1';
    layer0_outputs(2355) <= (inputs(87)) and not (inputs(206));
    layer0_outputs(2356) <= (inputs(36)) xor (inputs(129));
    layer0_outputs(2357) <= (inputs(4)) and not (inputs(135));
    layer0_outputs(2358) <= (inputs(51)) and not (inputs(44));
    layer0_outputs(2359) <= inputs(136);
    layer0_outputs(2360) <= not(inputs(8));
    layer0_outputs(2361) <= (inputs(77)) and not (inputs(128));
    layer0_outputs(2362) <= not((inputs(32)) xor (inputs(136)));
    layer0_outputs(2363) <= not(inputs(204));
    layer0_outputs(2364) <= not((inputs(8)) xor (inputs(23)));
    layer0_outputs(2365) <= (inputs(71)) or (inputs(242));
    layer0_outputs(2366) <= (inputs(78)) or (inputs(186));
    layer0_outputs(2367) <= not((inputs(45)) xor (inputs(69)));
    layer0_outputs(2368) <= (inputs(36)) or (inputs(95));
    layer0_outputs(2369) <= (inputs(16)) xor (inputs(115));
    layer0_outputs(2370) <= not(inputs(210));
    layer0_outputs(2371) <= (inputs(255)) or (inputs(53));
    layer0_outputs(2372) <= not(inputs(213)) or (inputs(143));
    layer0_outputs(2373) <= not(inputs(30)) or (inputs(186));
    layer0_outputs(2374) <= not((inputs(215)) or (inputs(80)));
    layer0_outputs(2375) <= not((inputs(50)) and (inputs(206)));
    layer0_outputs(2376) <= (inputs(180)) or (inputs(179));
    layer0_outputs(2377) <= not((inputs(127)) xor (inputs(11)));
    layer0_outputs(2378) <= (inputs(79)) or (inputs(135));
    layer0_outputs(2379) <= (inputs(20)) xor (inputs(127));
    layer0_outputs(2380) <= not((inputs(52)) or (inputs(229)));
    layer0_outputs(2381) <= not((inputs(106)) or (inputs(108)));
    layer0_outputs(2382) <= inputs(139);
    layer0_outputs(2383) <= not(inputs(15)) or (inputs(65));
    layer0_outputs(2384) <= (inputs(91)) or (inputs(99));
    layer0_outputs(2385) <= (inputs(246)) or (inputs(84));
    layer0_outputs(2386) <= not((inputs(224)) xor (inputs(135)));
    layer0_outputs(2387) <= not((inputs(221)) xor (inputs(166)));
    layer0_outputs(2388) <= (inputs(72)) xor (inputs(211));
    layer0_outputs(2389) <= not((inputs(227)) xor (inputs(171)));
    layer0_outputs(2390) <= inputs(118);
    layer0_outputs(2391) <= inputs(108);
    layer0_outputs(2392) <= (inputs(161)) or (inputs(229));
    layer0_outputs(2393) <= inputs(134);
    layer0_outputs(2394) <= not((inputs(58)) or (inputs(213)));
    layer0_outputs(2395) <= inputs(204);
    layer0_outputs(2396) <= not(inputs(76));
    layer0_outputs(2397) <= not((inputs(145)) xor (inputs(205)));
    layer0_outputs(2398) <= (inputs(189)) xor (inputs(31));
    layer0_outputs(2399) <= inputs(8);
    layer0_outputs(2400) <= (inputs(24)) and not (inputs(206));
    layer0_outputs(2401) <= (inputs(88)) xor (inputs(39));
    layer0_outputs(2402) <= not((inputs(59)) or (inputs(170)));
    layer0_outputs(2403) <= not((inputs(148)) xor (inputs(252)));
    layer0_outputs(2404) <= (inputs(127)) and (inputs(167));
    layer0_outputs(2405) <= not(inputs(107)) or (inputs(21));
    layer0_outputs(2406) <= (inputs(30)) and not (inputs(230));
    layer0_outputs(2407) <= not((inputs(38)) or (inputs(52)));
    layer0_outputs(2408) <= '1';
    layer0_outputs(2409) <= inputs(178);
    layer0_outputs(2410) <= '0';
    layer0_outputs(2411) <= not(inputs(144)) or (inputs(81));
    layer0_outputs(2412) <= (inputs(26)) and not (inputs(223));
    layer0_outputs(2413) <= (inputs(143)) and not (inputs(101));
    layer0_outputs(2414) <= not(inputs(32)) or (inputs(23));
    layer0_outputs(2415) <= not((inputs(226)) xor (inputs(243)));
    layer0_outputs(2416) <= not((inputs(215)) or (inputs(75)));
    layer0_outputs(2417) <= not((inputs(75)) xor (inputs(159)));
    layer0_outputs(2418) <= inputs(80);
    layer0_outputs(2419) <= (inputs(206)) or (inputs(169));
    layer0_outputs(2420) <= not((inputs(242)) xor (inputs(85)));
    layer0_outputs(2421) <= not(inputs(71)) or (inputs(12));
    layer0_outputs(2422) <= (inputs(145)) and not (inputs(35));
    layer0_outputs(2423) <= (inputs(241)) or (inputs(73));
    layer0_outputs(2424) <= (inputs(187)) or (inputs(41));
    layer0_outputs(2425) <= not((inputs(136)) or (inputs(208)));
    layer0_outputs(2426) <= not(inputs(237));
    layer0_outputs(2427) <= inputs(98);
    layer0_outputs(2428) <= not((inputs(251)) xor (inputs(89)));
    layer0_outputs(2429) <= (inputs(25)) or (inputs(162));
    layer0_outputs(2430) <= not(inputs(43)) or (inputs(243));
    layer0_outputs(2431) <= (inputs(49)) xor (inputs(155));
    layer0_outputs(2432) <= (inputs(249)) or (inputs(87));
    layer0_outputs(2433) <= inputs(33);
    layer0_outputs(2434) <= not((inputs(90)) or (inputs(38)));
    layer0_outputs(2435) <= (inputs(77)) xor (inputs(129));
    layer0_outputs(2436) <= (inputs(93)) or (inputs(116));
    layer0_outputs(2437) <= (inputs(204)) or (inputs(27));
    layer0_outputs(2438) <= not(inputs(50));
    layer0_outputs(2439) <= not(inputs(158));
    layer0_outputs(2440) <= inputs(104);
    layer0_outputs(2441) <= (inputs(203)) or (inputs(249));
    layer0_outputs(2442) <= not(inputs(7));
    layer0_outputs(2443) <= not(inputs(165)) or (inputs(191));
    layer0_outputs(2444) <= not(inputs(148));
    layer0_outputs(2445) <= (inputs(86)) xor (inputs(18));
    layer0_outputs(2446) <= (inputs(88)) or (inputs(235));
    layer0_outputs(2447) <= not(inputs(116)) or (inputs(143));
    layer0_outputs(2448) <= not((inputs(155)) or (inputs(178)));
    layer0_outputs(2449) <= (inputs(73)) xor (inputs(128));
    layer0_outputs(2450) <= inputs(252);
    layer0_outputs(2451) <= (inputs(201)) and not (inputs(125));
    layer0_outputs(2452) <= not((inputs(169)) xor (inputs(167)));
    layer0_outputs(2453) <= (inputs(137)) and not (inputs(111));
    layer0_outputs(2454) <= not(inputs(197)) or (inputs(14));
    layer0_outputs(2455) <= (inputs(156)) or (inputs(173));
    layer0_outputs(2456) <= not((inputs(148)) or (inputs(219)));
    layer0_outputs(2457) <= not((inputs(46)) and (inputs(5)));
    layer0_outputs(2458) <= (inputs(228)) xor (inputs(140));
    layer0_outputs(2459) <= inputs(37);
    layer0_outputs(2460) <= (inputs(38)) and (inputs(118));
    layer0_outputs(2461) <= not((inputs(3)) or (inputs(134)));
    layer0_outputs(2462) <= not(inputs(63)) or (inputs(0));
    layer0_outputs(2463) <= (inputs(168)) and not (inputs(194));
    layer0_outputs(2464) <= not(inputs(132)) or (inputs(135));
    layer0_outputs(2465) <= not(inputs(181)) or (inputs(231));
    layer0_outputs(2466) <= (inputs(163)) and not (inputs(6));
    layer0_outputs(2467) <= not((inputs(1)) xor (inputs(124)));
    layer0_outputs(2468) <= not((inputs(11)) and (inputs(191)));
    layer0_outputs(2469) <= inputs(92);
    layer0_outputs(2470) <= not(inputs(248)) or (inputs(111));
    layer0_outputs(2471) <= not(inputs(121)) or (inputs(211));
    layer0_outputs(2472) <= (inputs(164)) xor (inputs(181));
    layer0_outputs(2473) <= inputs(138);
    layer0_outputs(2474) <= not(inputs(87)) or (inputs(206));
    layer0_outputs(2475) <= (inputs(70)) and not (inputs(218));
    layer0_outputs(2476) <= (inputs(3)) xor (inputs(100));
    layer0_outputs(2477) <= (inputs(166)) or (inputs(53));
    layer0_outputs(2478) <= not(inputs(155));
    layer0_outputs(2479) <= (inputs(38)) xor (inputs(209));
    layer0_outputs(2480) <= not((inputs(70)) xor (inputs(141)));
    layer0_outputs(2481) <= inputs(212);
    layer0_outputs(2482) <= inputs(118);
    layer0_outputs(2483) <= (inputs(231)) xor (inputs(63));
    layer0_outputs(2484) <= not((inputs(228)) or (inputs(41)));
    layer0_outputs(2485) <= not((inputs(3)) xor (inputs(251)));
    layer0_outputs(2486) <= not(inputs(179)) or (inputs(15));
    layer0_outputs(2487) <= (inputs(119)) and not (inputs(127));
    layer0_outputs(2488) <= not((inputs(175)) xor (inputs(37)));
    layer0_outputs(2489) <= (inputs(64)) or (inputs(107));
    layer0_outputs(2490) <= not((inputs(131)) or (inputs(119)));
    layer0_outputs(2491) <= (inputs(104)) or (inputs(158));
    layer0_outputs(2492) <= not((inputs(30)) xor (inputs(13)));
    layer0_outputs(2493) <= (inputs(131)) and not (inputs(176));
    layer0_outputs(2494) <= not(inputs(134)) or (inputs(12));
    layer0_outputs(2495) <= (inputs(227)) xor (inputs(231));
    layer0_outputs(2496) <= (inputs(39)) or (inputs(10));
    layer0_outputs(2497) <= not((inputs(53)) or (inputs(210)));
    layer0_outputs(2498) <= (inputs(88)) and not (inputs(94));
    layer0_outputs(2499) <= not((inputs(206)) or (inputs(180)));
    layer0_outputs(2500) <= not(inputs(89));
    layer0_outputs(2501) <= inputs(213);
    layer0_outputs(2502) <= (inputs(127)) or (inputs(122));
    layer0_outputs(2503) <= not(inputs(118));
    layer0_outputs(2504) <= not(inputs(128));
    layer0_outputs(2505) <= not((inputs(102)) xor (inputs(192)));
    layer0_outputs(2506) <= not(inputs(126));
    layer0_outputs(2507) <= not(inputs(166)) or (inputs(229));
    layer0_outputs(2508) <= not(inputs(101)) or (inputs(198));
    layer0_outputs(2509) <= (inputs(225)) or (inputs(120));
    layer0_outputs(2510) <= inputs(107);
    layer0_outputs(2511) <= not(inputs(127)) or (inputs(7));
    layer0_outputs(2512) <= (inputs(184)) and not (inputs(2));
    layer0_outputs(2513) <= not(inputs(199)) or (inputs(192));
    layer0_outputs(2514) <= (inputs(234)) and (inputs(226));
    layer0_outputs(2515) <= inputs(142);
    layer0_outputs(2516) <= not(inputs(214)) or (inputs(24));
    layer0_outputs(2517) <= inputs(61);
    layer0_outputs(2518) <= (inputs(48)) or (inputs(0));
    layer0_outputs(2519) <= (inputs(102)) and not (inputs(161));
    layer0_outputs(2520) <= not(inputs(44));
    layer0_outputs(2521) <= (inputs(91)) and not (inputs(17));
    layer0_outputs(2522) <= (inputs(55)) or (inputs(239));
    layer0_outputs(2523) <= not(inputs(77)) or (inputs(202));
    layer0_outputs(2524) <= (inputs(143)) and (inputs(35));
    layer0_outputs(2525) <= (inputs(86)) or (inputs(229));
    layer0_outputs(2526) <= (inputs(217)) and not (inputs(51));
    layer0_outputs(2527) <= not(inputs(38));
    layer0_outputs(2528) <= not((inputs(171)) or (inputs(232)));
    layer0_outputs(2529) <= inputs(119);
    layer0_outputs(2530) <= not(inputs(198));
    layer0_outputs(2531) <= (inputs(206)) and (inputs(10));
    layer0_outputs(2532) <= (inputs(114)) xor (inputs(210));
    layer0_outputs(2533) <= inputs(49);
    layer0_outputs(2534) <= not(inputs(118)) or (inputs(99));
    layer0_outputs(2535) <= not(inputs(103));
    layer0_outputs(2536) <= not(inputs(165)) or (inputs(30));
    layer0_outputs(2537) <= (inputs(216)) or (inputs(208));
    layer0_outputs(2538) <= not((inputs(58)) or (inputs(110)));
    layer0_outputs(2539) <= not(inputs(168));
    layer0_outputs(2540) <= not((inputs(213)) or (inputs(227)));
    layer0_outputs(2541) <= (inputs(234)) xor (inputs(110));
    layer0_outputs(2542) <= '1';
    layer0_outputs(2543) <= (inputs(119)) and not (inputs(97));
    layer0_outputs(2544) <= (inputs(170)) and not (inputs(60));
    layer0_outputs(2545) <= (inputs(171)) or (inputs(144));
    layer0_outputs(2546) <= inputs(40);
    layer0_outputs(2547) <= not(inputs(219)) or (inputs(12));
    layer0_outputs(2548) <= (inputs(166)) and not (inputs(106));
    layer0_outputs(2549) <= (inputs(211)) or (inputs(170));
    layer0_outputs(2550) <= not(inputs(232));
    layer0_outputs(2551) <= (inputs(239)) and not (inputs(1));
    layer0_outputs(2552) <= inputs(129);
    layer0_outputs(2553) <= not(inputs(133)) or (inputs(173));
    layer0_outputs(2554) <= not((inputs(30)) and (inputs(14)));
    layer0_outputs(2555) <= inputs(192);
    layer0_outputs(2556) <= not((inputs(8)) or (inputs(186)));
    layer0_outputs(2557) <= not(inputs(168)) or (inputs(110));
    layer0_outputs(2558) <= (inputs(195)) and not (inputs(246));
    layer0_outputs(2559) <= (inputs(230)) and not (inputs(176));
    outputs(0) <= not(layer0_outputs(1783));
    outputs(1) <= layer0_outputs(462);
    outputs(2) <= (layer0_outputs(206)) xor (layer0_outputs(595));
    outputs(3) <= layer0_outputs(211);
    outputs(4) <= not(layer0_outputs(2033)) or (layer0_outputs(2044));
    outputs(5) <= not((layer0_outputs(408)) or (layer0_outputs(1577)));
    outputs(6) <= layer0_outputs(1491);
    outputs(7) <= not(layer0_outputs(1475));
    outputs(8) <= not((layer0_outputs(2487)) or (layer0_outputs(872)));
    outputs(9) <= not((layer0_outputs(1595)) or (layer0_outputs(2302)));
    outputs(10) <= (layer0_outputs(1733)) and not (layer0_outputs(61));
    outputs(11) <= not(layer0_outputs(1843));
    outputs(12) <= not((layer0_outputs(334)) or (layer0_outputs(2460)));
    outputs(13) <= not(layer0_outputs(598));
    outputs(14) <= (layer0_outputs(1245)) and not (layer0_outputs(1585));
    outputs(15) <= not(layer0_outputs(1607));
    outputs(16) <= not(layer0_outputs(2397)) or (layer0_outputs(1009));
    outputs(17) <= layer0_outputs(2294);
    outputs(18) <= (layer0_outputs(2091)) xor (layer0_outputs(2216));
    outputs(19) <= not(layer0_outputs(2403));
    outputs(20) <= (layer0_outputs(1088)) xor (layer0_outputs(2527));
    outputs(21) <= not(layer0_outputs(2004));
    outputs(22) <= layer0_outputs(1461);
    outputs(23) <= (layer0_outputs(284)) xor (layer0_outputs(1997));
    outputs(24) <= not(layer0_outputs(263));
    outputs(25) <= layer0_outputs(541);
    outputs(26) <= (layer0_outputs(1248)) or (layer0_outputs(1291));
    outputs(27) <= layer0_outputs(2336);
    outputs(28) <= not((layer0_outputs(754)) or (layer0_outputs(585)));
    outputs(29) <= (layer0_outputs(1563)) or (layer0_outputs(2399));
    outputs(30) <= not(layer0_outputs(129)) or (layer0_outputs(81));
    outputs(31) <= not(layer0_outputs(2042)) or (layer0_outputs(676));
    outputs(32) <= not(layer0_outputs(2444));
    outputs(33) <= not((layer0_outputs(127)) and (layer0_outputs(597)));
    outputs(34) <= layer0_outputs(1001);
    outputs(35) <= not(layer0_outputs(492)) or (layer0_outputs(1255));
    outputs(36) <= not(layer0_outputs(2137));
    outputs(37) <= not((layer0_outputs(2171)) and (layer0_outputs(1123)));
    outputs(38) <= not(layer0_outputs(1514));
    outputs(39) <= (layer0_outputs(1573)) or (layer0_outputs(1687));
    outputs(40) <= not(layer0_outputs(1185)) or (layer0_outputs(431));
    outputs(41) <= layer0_outputs(1699);
    outputs(42) <= (layer0_outputs(751)) and (layer0_outputs(994));
    outputs(43) <= not(layer0_outputs(168));
    outputs(44) <= layer0_outputs(1500);
    outputs(45) <= not(layer0_outputs(1724));
    outputs(46) <= not(layer0_outputs(384));
    outputs(47) <= not(layer0_outputs(1987)) or (layer0_outputs(1432));
    outputs(48) <= (layer0_outputs(1112)) and not (layer0_outputs(716));
    outputs(49) <= layer0_outputs(1096);
    outputs(50) <= not((layer0_outputs(1679)) and (layer0_outputs(1057)));
    outputs(51) <= not(layer0_outputs(319)) or (layer0_outputs(500));
    outputs(52) <= not(layer0_outputs(1786));
    outputs(53) <= not(layer0_outputs(279)) or (layer0_outputs(602));
    outputs(54) <= (layer0_outputs(2556)) xor (layer0_outputs(2520));
    outputs(55) <= not(layer0_outputs(272));
    outputs(56) <= (layer0_outputs(457)) and not (layer0_outputs(2272));
    outputs(57) <= (layer0_outputs(846)) and not (layer0_outputs(273));
    outputs(58) <= layer0_outputs(320);
    outputs(59) <= layer0_outputs(134);
    outputs(60) <= layer0_outputs(793);
    outputs(61) <= layer0_outputs(1144);
    outputs(62) <= (layer0_outputs(433)) xor (layer0_outputs(48));
    outputs(63) <= not(layer0_outputs(1783)) or (layer0_outputs(1604));
    outputs(64) <= not(layer0_outputs(1751));
    outputs(65) <= not(layer0_outputs(2491)) or (layer0_outputs(632));
    outputs(66) <= not((layer0_outputs(1374)) xor (layer0_outputs(1106)));
    outputs(67) <= not(layer0_outputs(1967)) or (layer0_outputs(2276));
    outputs(68) <= (layer0_outputs(2311)) and not (layer0_outputs(2099));
    outputs(69) <= not((layer0_outputs(1559)) and (layer0_outputs(629)));
    outputs(70) <= (layer0_outputs(1981)) or (layer0_outputs(1883));
    outputs(71) <= not(layer0_outputs(550)) or (layer0_outputs(1070));
    outputs(72) <= not(layer0_outputs(2257));
    outputs(73) <= not((layer0_outputs(2093)) xor (layer0_outputs(1400)));
    outputs(74) <= not(layer0_outputs(593));
    outputs(75) <= layer0_outputs(671);
    outputs(76) <= not(layer0_outputs(2163));
    outputs(77) <= layer0_outputs(1515);
    outputs(78) <= (layer0_outputs(2025)) and not (layer0_outputs(565));
    outputs(79) <= (layer0_outputs(2140)) or (layer0_outputs(901));
    outputs(80) <= not((layer0_outputs(2397)) xor (layer0_outputs(846)));
    outputs(81) <= (layer0_outputs(2225)) or (layer0_outputs(1179));
    outputs(82) <= layer0_outputs(282);
    outputs(83) <= (layer0_outputs(1111)) or (layer0_outputs(1130));
    outputs(84) <= not(layer0_outputs(2046));
    outputs(85) <= not(layer0_outputs(1140));
    outputs(86) <= (layer0_outputs(479)) and not (layer0_outputs(1525));
    outputs(87) <= not(layer0_outputs(242));
    outputs(88) <= (layer0_outputs(1883)) xor (layer0_outputs(911));
    outputs(89) <= (layer0_outputs(1778)) and not (layer0_outputs(1072));
    outputs(90) <= not((layer0_outputs(251)) xor (layer0_outputs(1753)));
    outputs(91) <= not((layer0_outputs(802)) and (layer0_outputs(2141)));
    outputs(92) <= layer0_outputs(1205);
    outputs(93) <= not(layer0_outputs(432));
    outputs(94) <= (layer0_outputs(1488)) and not (layer0_outputs(845));
    outputs(95) <= not(layer0_outputs(1197)) or (layer0_outputs(1269));
    outputs(96) <= not(layer0_outputs(517));
    outputs(97) <= not((layer0_outputs(612)) xor (layer0_outputs(2324)));
    outputs(98) <= not(layer0_outputs(2111));
    outputs(99) <= not((layer0_outputs(419)) and (layer0_outputs(2516)));
    outputs(100) <= (layer0_outputs(571)) xor (layer0_outputs(581));
    outputs(101) <= layer0_outputs(974);
    outputs(102) <= not((layer0_outputs(1377)) or (layer0_outputs(1425)));
    outputs(103) <= (layer0_outputs(1185)) xor (layer0_outputs(2));
    outputs(104) <= not(layer0_outputs(2464));
    outputs(105) <= not((layer0_outputs(1897)) xor (layer0_outputs(1670)));
    outputs(106) <= layer0_outputs(1238);
    outputs(107) <= (layer0_outputs(764)) and not (layer0_outputs(1007));
    outputs(108) <= layer0_outputs(926);
    outputs(109) <= layer0_outputs(2152);
    outputs(110) <= not(layer0_outputs(165));
    outputs(111) <= (layer0_outputs(2545)) xor (layer0_outputs(1039));
    outputs(112) <= (layer0_outputs(1203)) and not (layer0_outputs(1864));
    outputs(113) <= not(layer0_outputs(383));
    outputs(114) <= not(layer0_outputs(2502));
    outputs(115) <= layer0_outputs(2382);
    outputs(116) <= not((layer0_outputs(994)) xor (layer0_outputs(760)));
    outputs(117) <= layer0_outputs(2075);
    outputs(118) <= (layer0_outputs(1141)) and (layer0_outputs(1983));
    outputs(119) <= layer0_outputs(2044);
    outputs(120) <= not(layer0_outputs(1802));
    outputs(121) <= (layer0_outputs(2355)) and not (layer0_outputs(2178));
    outputs(122) <= not(layer0_outputs(1242));
    outputs(123) <= not((layer0_outputs(1127)) xor (layer0_outputs(220)));
    outputs(124) <= not(layer0_outputs(321)) or (layer0_outputs(1110));
    outputs(125) <= layer0_outputs(27);
    outputs(126) <= not((layer0_outputs(2235)) xor (layer0_outputs(1214)));
    outputs(127) <= (layer0_outputs(1306)) xor (layer0_outputs(1585));
    outputs(128) <= (layer0_outputs(1780)) and not (layer0_outputs(260));
    outputs(129) <= not((layer0_outputs(324)) xor (layer0_outputs(1601)));
    outputs(130) <= not((layer0_outputs(2078)) xor (layer0_outputs(1214)));
    outputs(131) <= not((layer0_outputs(472)) xor (layer0_outputs(1592)));
    outputs(132) <= (layer0_outputs(2497)) or (layer0_outputs(31));
    outputs(133) <= not((layer0_outputs(1605)) or (layer0_outputs(1022)));
    outputs(134) <= (layer0_outputs(1972)) and not (layer0_outputs(2258));
    outputs(135) <= not(layer0_outputs(1938)) or (layer0_outputs(1301));
    outputs(136) <= not(layer0_outputs(1951));
    outputs(137) <= not((layer0_outputs(1861)) or (layer0_outputs(1770)));
    outputs(138) <= not(layer0_outputs(870));
    outputs(139) <= not((layer0_outputs(466)) xor (layer0_outputs(725)));
    outputs(140) <= not(layer0_outputs(1021)) or (layer0_outputs(2244));
    outputs(141) <= not(layer0_outputs(139));
    outputs(142) <= layer0_outputs(1870);
    outputs(143) <= layer0_outputs(2376);
    outputs(144) <= layer0_outputs(499);
    outputs(145) <= layer0_outputs(2223);
    outputs(146) <= layer0_outputs(362);
    outputs(147) <= layer0_outputs(1742);
    outputs(148) <= not((layer0_outputs(1933)) or (layer0_outputs(1926)));
    outputs(149) <= not(layer0_outputs(1516)) or (layer0_outputs(2012));
    outputs(150) <= (layer0_outputs(1508)) or (layer0_outputs(769));
    outputs(151) <= not(layer0_outputs(2073));
    outputs(152) <= layer0_outputs(1387);
    outputs(153) <= layer0_outputs(1965);
    outputs(154) <= not(layer0_outputs(62));
    outputs(155) <= (layer0_outputs(134)) and not (layer0_outputs(605));
    outputs(156) <= layer0_outputs(234);
    outputs(157) <= (layer0_outputs(1846)) and not (layer0_outputs(61));
    outputs(158) <= (layer0_outputs(369)) and (layer0_outputs(1263));
    outputs(159) <= not(layer0_outputs(601));
    outputs(160) <= not(layer0_outputs(599)) or (layer0_outputs(730));
    outputs(161) <= not(layer0_outputs(255));
    outputs(162) <= layer0_outputs(1392);
    outputs(163) <= layer0_outputs(411);
    outputs(164) <= not(layer0_outputs(1998));
    outputs(165) <= (layer0_outputs(521)) and (layer0_outputs(954));
    outputs(166) <= not((layer0_outputs(9)) and (layer0_outputs(1490)));
    outputs(167) <= not(layer0_outputs(2028));
    outputs(168) <= not((layer0_outputs(220)) or (layer0_outputs(1417)));
    outputs(169) <= not(layer0_outputs(1056));
    outputs(170) <= not(layer0_outputs(1267));
    outputs(171) <= layer0_outputs(874);
    outputs(172) <= (layer0_outputs(385)) and not (layer0_outputs(2393));
    outputs(173) <= (layer0_outputs(1955)) and not (layer0_outputs(1514));
    outputs(174) <= layer0_outputs(583);
    outputs(175) <= layer0_outputs(2187);
    outputs(176) <= not(layer0_outputs(448)) or (layer0_outputs(1134));
    outputs(177) <= layer0_outputs(1513);
    outputs(178) <= not((layer0_outputs(1201)) or (layer0_outputs(1811)));
    outputs(179) <= not(layer0_outputs(892)) or (layer0_outputs(632));
    outputs(180) <= not(layer0_outputs(2188));
    outputs(181) <= layer0_outputs(1095);
    outputs(182) <= (layer0_outputs(143)) or (layer0_outputs(1513));
    outputs(183) <= (layer0_outputs(2527)) and not (layer0_outputs(105));
    outputs(184) <= not(layer0_outputs(1621));
    outputs(185) <= layer0_outputs(1070);
    outputs(186) <= not(layer0_outputs(1023));
    outputs(187) <= (layer0_outputs(596)) and not (layer0_outputs(311));
    outputs(188) <= not(layer0_outputs(975));
    outputs(189) <= not((layer0_outputs(1124)) xor (layer0_outputs(1235)));
    outputs(190) <= layer0_outputs(1466);
    outputs(191) <= not(layer0_outputs(2217));
    outputs(192) <= (layer0_outputs(842)) and not (layer0_outputs(104));
    outputs(193) <= (layer0_outputs(2539)) and not (layer0_outputs(1497));
    outputs(194) <= not(layer0_outputs(1775));
    outputs(195) <= not(layer0_outputs(1909)) or (layer0_outputs(1248));
    outputs(196) <= layer0_outputs(677);
    outputs(197) <= not(layer0_outputs(1472));
    outputs(198) <= (layer0_outputs(2126)) or (layer0_outputs(247));
    outputs(199) <= not((layer0_outputs(419)) and (layer0_outputs(353)));
    outputs(200) <= layer0_outputs(1959);
    outputs(201) <= (layer0_outputs(2321)) and not (layer0_outputs(946));
    outputs(202) <= layer0_outputs(986);
    outputs(203) <= not((layer0_outputs(366)) and (layer0_outputs(747)));
    outputs(204) <= layer0_outputs(1168);
    outputs(205) <= (layer0_outputs(1515)) and not (layer0_outputs(2159));
    outputs(206) <= layer0_outputs(470);
    outputs(207) <= not(layer0_outputs(2280));
    outputs(208) <= not(layer0_outputs(1087));
    outputs(209) <= (layer0_outputs(1489)) xor (layer0_outputs(1463));
    outputs(210) <= (layer0_outputs(1668)) and (layer0_outputs(270));
    outputs(211) <= not((layer0_outputs(1967)) and (layer0_outputs(1673)));
    outputs(212) <= (layer0_outputs(2407)) and not (layer0_outputs(512));
    outputs(213) <= (layer0_outputs(1227)) and (layer0_outputs(2156));
    outputs(214) <= (layer0_outputs(412)) and (layer0_outputs(552));
    outputs(215) <= (layer0_outputs(144)) xor (layer0_outputs(64));
    outputs(216) <= not(layer0_outputs(1836));
    outputs(217) <= layer0_outputs(2387);
    outputs(218) <= layer0_outputs(2350);
    outputs(219) <= not(layer0_outputs(2502));
    outputs(220) <= layer0_outputs(1357);
    outputs(221) <= (layer0_outputs(317)) and (layer0_outputs(190));
    outputs(222) <= not(layer0_outputs(2342));
    outputs(223) <= not(layer0_outputs(644));
    outputs(224) <= not(layer0_outputs(430)) or (layer0_outputs(293));
    outputs(225) <= not((layer0_outputs(1789)) xor (layer0_outputs(815)));
    outputs(226) <= not((layer0_outputs(939)) xor (layer0_outputs(1556)));
    outputs(227) <= not((layer0_outputs(730)) or (layer0_outputs(1047)));
    outputs(228) <= not(layer0_outputs(1623)) or (layer0_outputs(142));
    outputs(229) <= (layer0_outputs(468)) and not (layer0_outputs(697));
    outputs(230) <= (layer0_outputs(1509)) xor (layer0_outputs(2532));
    outputs(231) <= not((layer0_outputs(1520)) and (layer0_outputs(1963)));
    outputs(232) <= not(layer0_outputs(1451));
    outputs(233) <= (layer0_outputs(34)) or (layer0_outputs(2246));
    outputs(234) <= (layer0_outputs(724)) xor (layer0_outputs(1400));
    outputs(235) <= not((layer0_outputs(290)) xor (layer0_outputs(1161)));
    outputs(236) <= not((layer0_outputs(1075)) and (layer0_outputs(1443)));
    outputs(237) <= layer0_outputs(1082);
    outputs(238) <= (layer0_outputs(879)) and (layer0_outputs(1712));
    outputs(239) <= not(layer0_outputs(857));
    outputs(240) <= layer0_outputs(403);
    outputs(241) <= (layer0_outputs(615)) and (layer0_outputs(308));
    outputs(242) <= not(layer0_outputs(1302));
    outputs(243) <= (layer0_outputs(1502)) or (layer0_outputs(511));
    outputs(244) <= layer0_outputs(2390);
    outputs(245) <= (layer0_outputs(1307)) or (layer0_outputs(659));
    outputs(246) <= (layer0_outputs(2455)) and not (layer0_outputs(2548));
    outputs(247) <= not(layer0_outputs(94));
    outputs(248) <= (layer0_outputs(536)) and (layer0_outputs(571));
    outputs(249) <= layer0_outputs(1452);
    outputs(250) <= not(layer0_outputs(1657)) or (layer0_outputs(528));
    outputs(251) <= not(layer0_outputs(2084));
    outputs(252) <= (layer0_outputs(1744)) and (layer0_outputs(554));
    outputs(253) <= not(layer0_outputs(107));
    outputs(254) <= layer0_outputs(464);
    outputs(255) <= not((layer0_outputs(2254)) xor (layer0_outputs(625)));
    outputs(256) <= (layer0_outputs(268)) and not (layer0_outputs(379));
    outputs(257) <= layer0_outputs(217);
    outputs(258) <= (layer0_outputs(2236)) and not (layer0_outputs(1262));
    outputs(259) <= (layer0_outputs(569)) xor (layer0_outputs(2330));
    outputs(260) <= not((layer0_outputs(2501)) xor (layer0_outputs(1575)));
    outputs(261) <= layer0_outputs(1801);
    outputs(262) <= not(layer0_outputs(940));
    outputs(263) <= (layer0_outputs(1381)) and not (layer0_outputs(1295));
    outputs(264) <= (layer0_outputs(1614)) or (layer0_outputs(1676));
    outputs(265) <= not((layer0_outputs(1772)) or (layer0_outputs(1015)));
    outputs(266) <= (layer0_outputs(1173)) and not (layer0_outputs(48));
    outputs(267) <= not((layer0_outputs(210)) or (layer0_outputs(2229)));
    outputs(268) <= not((layer0_outputs(888)) or (layer0_outputs(64)));
    outputs(269) <= not(layer0_outputs(95));
    outputs(270) <= not((layer0_outputs(45)) xor (layer0_outputs(2415)));
    outputs(271) <= not(layer0_outputs(1046));
    outputs(272) <= (layer0_outputs(2494)) and not (layer0_outputs(354));
    outputs(273) <= (layer0_outputs(262)) and (layer0_outputs(290));
    outputs(274) <= (layer0_outputs(2192)) and not (layer0_outputs(1011));
    outputs(275) <= not((layer0_outputs(2210)) xor (layer0_outputs(1777)));
    outputs(276) <= (layer0_outputs(1204)) xor (layer0_outputs(1439));
    outputs(277) <= (layer0_outputs(2162)) and not (layer0_outputs(1824));
    outputs(278) <= not(layer0_outputs(2295));
    outputs(279) <= not((layer0_outputs(1001)) xor (layer0_outputs(2124)));
    outputs(280) <= layer0_outputs(352);
    outputs(281) <= layer0_outputs(413);
    outputs(282) <= '0';
    outputs(283) <= (layer0_outputs(130)) and not (layer0_outputs(2433));
    outputs(284) <= (layer0_outputs(1996)) and (layer0_outputs(2195));
    outputs(285) <= not(layer0_outputs(2077));
    outputs(286) <= layer0_outputs(72);
    outputs(287) <= (layer0_outputs(838)) and (layer0_outputs(624));
    outputs(288) <= not(layer0_outputs(1848));
    outputs(289) <= not((layer0_outputs(1629)) or (layer0_outputs(501)));
    outputs(290) <= layer0_outputs(392);
    outputs(291) <= not((layer0_outputs(1062)) or (layer0_outputs(2293)));
    outputs(292) <= (layer0_outputs(2333)) and not (layer0_outputs(1013));
    outputs(293) <= layer0_outputs(2157);
    outputs(294) <= (layer0_outputs(818)) and not (layer0_outputs(310));
    outputs(295) <= (layer0_outputs(1761)) and not (layer0_outputs(160));
    outputs(296) <= (layer0_outputs(1764)) and (layer0_outputs(1334));
    outputs(297) <= (layer0_outputs(1645)) and not (layer0_outputs(1484));
    outputs(298) <= not((layer0_outputs(1158)) or (layer0_outputs(935)));
    outputs(299) <= not(layer0_outputs(88));
    outputs(300) <= not((layer0_outputs(2525)) or (layer0_outputs(2108)));
    outputs(301) <= not(layer0_outputs(1700));
    outputs(302) <= (layer0_outputs(873)) and (layer0_outputs(1608));
    outputs(303) <= not((layer0_outputs(300)) or (layer0_outputs(1869)));
    outputs(304) <= (layer0_outputs(1418)) and not (layer0_outputs(1060));
    outputs(305) <= (layer0_outputs(1439)) and not (layer0_outputs(296));
    outputs(306) <= (layer0_outputs(1906)) and not (layer0_outputs(1793));
    outputs(307) <= not((layer0_outputs(1798)) or (layer0_outputs(1463)));
    outputs(308) <= not((layer0_outputs(94)) xor (layer0_outputs(1819)));
    outputs(309) <= layer0_outputs(345);
    outputs(310) <= not(layer0_outputs(2476));
    outputs(311) <= not(layer0_outputs(666));
    outputs(312) <= (layer0_outputs(2151)) and not (layer0_outputs(399));
    outputs(313) <= not((layer0_outputs(596)) xor (layer0_outputs(1806)));
    outputs(314) <= not((layer0_outputs(148)) or (layer0_outputs(1527)));
    outputs(315) <= (layer0_outputs(2498)) and not (layer0_outputs(1202));
    outputs(316) <= (layer0_outputs(316)) and not (layer0_outputs(338));
    outputs(317) <= not(layer0_outputs(191));
    outputs(318) <= (layer0_outputs(1042)) and not (layer0_outputs(78));
    outputs(319) <= not((layer0_outputs(2038)) xor (layer0_outputs(1633)));
    outputs(320) <= (layer0_outputs(1705)) and not (layer0_outputs(30));
    outputs(321) <= (layer0_outputs(2103)) and not (layer0_outputs(89));
    outputs(322) <= (layer0_outputs(1769)) and (layer0_outputs(2136));
    outputs(323) <= (layer0_outputs(1568)) and (layer0_outputs(1566));
    outputs(324) <= layer0_outputs(1414);
    outputs(325) <= (layer0_outputs(259)) and (layer0_outputs(108));
    outputs(326) <= (layer0_outputs(782)) or (layer0_outputs(1119));
    outputs(327) <= (layer0_outputs(590)) and not (layer0_outputs(1934));
    outputs(328) <= (layer0_outputs(2081)) and not (layer0_outputs(277));
    outputs(329) <= (layer0_outputs(2155)) and not (layer0_outputs(542));
    outputs(330) <= not((layer0_outputs(768)) or (layer0_outputs(24)));
    outputs(331) <= (layer0_outputs(1873)) and not (layer0_outputs(2510));
    outputs(332) <= (layer0_outputs(543)) and not (layer0_outputs(2459));
    outputs(333) <= (layer0_outputs(2049)) and (layer0_outputs(509));
    outputs(334) <= not((layer0_outputs(2441)) or (layer0_outputs(955)));
    outputs(335) <= (layer0_outputs(1534)) and not (layer0_outputs(718));
    outputs(336) <= not((layer0_outputs(146)) or (layer0_outputs(1290)));
    outputs(337) <= (layer0_outputs(1369)) and not (layer0_outputs(2266));
    outputs(338) <= (layer0_outputs(1304)) and not (layer0_outputs(2290));
    outputs(339) <= (layer0_outputs(577)) and not (layer0_outputs(161));
    outputs(340) <= (layer0_outputs(1665)) and (layer0_outputs(1008));
    outputs(341) <= (layer0_outputs(2248)) xor (layer0_outputs(1754));
    outputs(342) <= not(layer0_outputs(237));
    outputs(343) <= not((layer0_outputs(1817)) or (layer0_outputs(147)));
    outputs(344) <= (layer0_outputs(534)) and not (layer0_outputs(2489));
    outputs(345) <= not((layer0_outputs(107)) or (layer0_outputs(2455)));
    outputs(346) <= not(layer0_outputs(1914));
    outputs(347) <= (layer0_outputs(1377)) and not (layer0_outputs(1011));
    outputs(348) <= not((layer0_outputs(179)) or (layer0_outputs(677)));
    outputs(349) <= (layer0_outputs(2514)) and not (layer0_outputs(289));
    outputs(350) <= not(layer0_outputs(1139));
    outputs(351) <= (layer0_outputs(381)) and not (layer0_outputs(1183));
    outputs(352) <= (layer0_outputs(1344)) and not (layer0_outputs(1818));
    outputs(353) <= (layer0_outputs(232)) and not (layer0_outputs(375));
    outputs(354) <= (layer0_outputs(1902)) and not (layer0_outputs(1188));
    outputs(355) <= (layer0_outputs(1310)) and not (layer0_outputs(1287));
    outputs(356) <= (layer0_outputs(945)) and not (layer0_outputs(2288));
    outputs(357) <= layer0_outputs(1792);
    outputs(358) <= not((layer0_outputs(1923)) xor (layer0_outputs(1505)));
    outputs(359) <= layer0_outputs(1933);
    outputs(360) <= (layer0_outputs(2192)) and not (layer0_outputs(277));
    outputs(361) <= (layer0_outputs(932)) and (layer0_outputs(394));
    outputs(362) <= (layer0_outputs(1830)) and not (layer0_outputs(694));
    outputs(363) <= '0';
    outputs(364) <= not((layer0_outputs(161)) or (layer0_outputs(415)));
    outputs(365) <= not((layer0_outputs(1285)) xor (layer0_outputs(573)));
    outputs(366) <= not((layer0_outputs(56)) or (layer0_outputs(1024)));
    outputs(367) <= not(layer0_outputs(2453));
    outputs(368) <= (layer0_outputs(1441)) and not (layer0_outputs(6));
    outputs(369) <= not((layer0_outputs(1501)) or (layer0_outputs(959)));
    outputs(370) <= not((layer0_outputs(1934)) or (layer0_outputs(2034)));
    outputs(371) <= not(layer0_outputs(675));
    outputs(372) <= not((layer0_outputs(2139)) xor (layer0_outputs(1702)));
    outputs(373) <= not((layer0_outputs(461)) or (layer0_outputs(2057)));
    outputs(374) <= (layer0_outputs(2082)) and (layer0_outputs(1717));
    outputs(375) <= layer0_outputs(185);
    outputs(376) <= (layer0_outputs(2214)) and (layer0_outputs(391));
    outputs(377) <= (layer0_outputs(2113)) and not (layer0_outputs(266));
    outputs(378) <= not(layer0_outputs(1080));
    outputs(379) <= not(layer0_outputs(370));
    outputs(380) <= (layer0_outputs(2112)) and (layer0_outputs(2405));
    outputs(381) <= layer0_outputs(1863);
    outputs(382) <= not((layer0_outputs(1038)) or (layer0_outputs(399)));
    outputs(383) <= (layer0_outputs(1723)) and not (layer0_outputs(343));
    outputs(384) <= (layer0_outputs(1520)) and (layer0_outputs(1299));
    outputs(385) <= not((layer0_outputs(1501)) or (layer0_outputs(81)));
    outputs(386) <= (layer0_outputs(1682)) and not (layer0_outputs(115));
    outputs(387) <= not((layer0_outputs(1949)) or (layer0_outputs(1353)));
    outputs(388) <= (layer0_outputs(2394)) and not (layer0_outputs(242));
    outputs(389) <= (layer0_outputs(870)) and not (layer0_outputs(285));
    outputs(390) <= not((layer0_outputs(816)) or (layer0_outputs(1847)));
    outputs(391) <= layer0_outputs(1149);
    outputs(392) <= (layer0_outputs(1086)) and (layer0_outputs(842));
    outputs(393) <= (layer0_outputs(2016)) and (layer0_outputs(2111));
    outputs(394) <= (layer0_outputs(2470)) and (layer0_outputs(2480));
    outputs(395) <= not((layer0_outputs(1960)) or (layer0_outputs(888)));
    outputs(396) <= (layer0_outputs(2416)) and (layer0_outputs(836));
    outputs(397) <= (layer0_outputs(232)) and (layer0_outputs(130));
    outputs(398) <= (layer0_outputs(427)) and not (layer0_outputs(1166));
    outputs(399) <= layer0_outputs(1606);
    outputs(400) <= (layer0_outputs(1996)) and not (layer0_outputs(700));
    outputs(401) <= not((layer0_outputs(455)) or (layer0_outputs(701)));
    outputs(402) <= layer0_outputs(2536);
    outputs(403) <= (layer0_outputs(474)) and (layer0_outputs(1270));
    outputs(404) <= (layer0_outputs(754)) and not (layer0_outputs(1461));
    outputs(405) <= (layer0_outputs(1225)) and not (layer0_outputs(1105));
    outputs(406) <= (layer0_outputs(885)) and not (layer0_outputs(1045));
    outputs(407) <= (layer0_outputs(804)) and not (layer0_outputs(1528));
    outputs(408) <= (layer0_outputs(2028)) and not (layer0_outputs(1728));
    outputs(409) <= not((layer0_outputs(410)) or (layer0_outputs(1116)));
    outputs(410) <= layer0_outputs(243);
    outputs(411) <= (layer0_outputs(2414)) xor (layer0_outputs(895));
    outputs(412) <= (layer0_outputs(423)) and not (layer0_outputs(1004));
    outputs(413) <= not((layer0_outputs(537)) xor (layer0_outputs(1857)));
    outputs(414) <= not((layer0_outputs(1874)) xor (layer0_outputs(1522)));
    outputs(415) <= not((layer0_outputs(565)) or (layer0_outputs(504)));
    outputs(416) <= layer0_outputs(2440);
    outputs(417) <= (layer0_outputs(745)) and (layer0_outputs(1908));
    outputs(418) <= (layer0_outputs(1541)) xor (layer0_outputs(2557));
    outputs(419) <= (layer0_outputs(1253)) and not (layer0_outputs(1551));
    outputs(420) <= (layer0_outputs(1724)) and not (layer0_outputs(378));
    outputs(421) <= (layer0_outputs(1970)) and not (layer0_outputs(477));
    outputs(422) <= (layer0_outputs(297)) and not (layer0_outputs(174));
    outputs(423) <= not(layer0_outputs(1663));
    outputs(424) <= (layer0_outputs(2134)) and not (layer0_outputs(2517));
    outputs(425) <= layer0_outputs(209);
    outputs(426) <= (layer0_outputs(2212)) and not (layer0_outputs(1721));
    outputs(427) <= not(layer0_outputs(1195));
    outputs(428) <= (layer0_outputs(1117)) and not (layer0_outputs(281));
    outputs(429) <= not((layer0_outputs(354)) or (layer0_outputs(387)));
    outputs(430) <= layer0_outputs(1006);
    outputs(431) <= (layer0_outputs(755)) and (layer0_outputs(1344));
    outputs(432) <= (layer0_outputs(985)) and not (layer0_outputs(664));
    outputs(433) <= not((layer0_outputs(1052)) or (layer0_outputs(1459)));
    outputs(434) <= not(layer0_outputs(2453));
    outputs(435) <= '0';
    outputs(436) <= not(layer0_outputs(2336));
    outputs(437) <= (layer0_outputs(1311)) and not (layer0_outputs(1617));
    outputs(438) <= (layer0_outputs(549)) and (layer0_outputs(145));
    outputs(439) <= (layer0_outputs(1862)) and not (layer0_outputs(1019));
    outputs(440) <= (layer0_outputs(506)) and not (layer0_outputs(1020));
    outputs(441) <= not((layer0_outputs(2035)) or (layer0_outputs(230)));
    outputs(442) <= not((layer0_outputs(527)) or (layer0_outputs(1062)));
    outputs(443) <= (layer0_outputs(1258)) and not (layer0_outputs(1727));
    outputs(444) <= (layer0_outputs(1160)) and not (layer0_outputs(437));
    outputs(445) <= layer0_outputs(535);
    outputs(446) <= (layer0_outputs(877)) and not (layer0_outputs(2495));
    outputs(447) <= (layer0_outputs(438)) and not (layer0_outputs(378));
    outputs(448) <= (layer0_outputs(1756)) xor (layer0_outputs(17));
    outputs(449) <= not((layer0_outputs(1701)) or (layer0_outputs(1151)));
    outputs(450) <= '0';
    outputs(451) <= not((layer0_outputs(1801)) xor (layer0_outputs(2087)));
    outputs(452) <= not((layer0_outputs(103)) or (layer0_outputs(11)));
    outputs(453) <= not((layer0_outputs(1808)) or (layer0_outputs(1321)));
    outputs(454) <= layer0_outputs(1775);
    outputs(455) <= not(layer0_outputs(1838));
    outputs(456) <= (layer0_outputs(1784)) xor (layer0_outputs(2103));
    outputs(457) <= (layer0_outputs(2516)) and not (layer0_outputs(1675));
    outputs(458) <= layer0_outputs(349);
    outputs(459) <= (layer0_outputs(1303)) and (layer0_outputs(532));
    outputs(460) <= (layer0_outputs(1759)) and not (layer0_outputs(2203));
    outputs(461) <= not((layer0_outputs(1649)) xor (layer0_outputs(1577)));
    outputs(462) <= not((layer0_outputs(1853)) or (layer0_outputs(2339)));
    outputs(463) <= (layer0_outputs(315)) and not (layer0_outputs(2428));
    outputs(464) <= not((layer0_outputs(1327)) and (layer0_outputs(2554)));
    outputs(465) <= not(layer0_outputs(1603));
    outputs(466) <= not((layer0_outputs(536)) xor (layer0_outputs(534)));
    outputs(467) <= (layer0_outputs(2059)) and not (layer0_outputs(989));
    outputs(468) <= (layer0_outputs(1199)) and (layer0_outputs(1315));
    outputs(469) <= not((layer0_outputs(1066)) or (layer0_outputs(1672)));
    outputs(470) <= '0';
    outputs(471) <= (layer0_outputs(2188)) and (layer0_outputs(75));
    outputs(472) <= (layer0_outputs(388)) and not (layer0_outputs(1275));
    outputs(473) <= (layer0_outputs(170)) and not (layer0_outputs(54));
    outputs(474) <= not((layer0_outputs(2190)) or (layer0_outputs(1468)));
    outputs(475) <= layer0_outputs(1882);
    outputs(476) <= layer0_outputs(122);
    outputs(477) <= not((layer0_outputs(1679)) or (layer0_outputs(2175)));
    outputs(478) <= (layer0_outputs(106)) and not (layer0_outputs(875));
    outputs(479) <= not(layer0_outputs(365));
    outputs(480) <= (layer0_outputs(771)) and (layer0_outputs(1689));
    outputs(481) <= not(layer0_outputs(494));
    outputs(482) <= not(layer0_outputs(1273));
    outputs(483) <= (layer0_outputs(5)) and not (layer0_outputs(193));
    outputs(484) <= (layer0_outputs(169)) and not (layer0_outputs(2559));
    outputs(485) <= not((layer0_outputs(1128)) xor (layer0_outputs(2250)));
    outputs(486) <= layer0_outputs(1337);
    outputs(487) <= (layer0_outputs(1531)) and not (layer0_outputs(377));
    outputs(488) <= (layer0_outputs(2421)) and not (layer0_outputs(1964));
    outputs(489) <= (layer0_outputs(257)) and not (layer0_outputs(919));
    outputs(490) <= (layer0_outputs(1251)) and not (layer0_outputs(1973));
    outputs(491) <= (layer0_outputs(2253)) and not (layer0_outputs(460));
    outputs(492) <= not(layer0_outputs(1465));
    outputs(493) <= (layer0_outputs(254)) and not (layer0_outputs(699));
    outputs(494) <= not((layer0_outputs(264)) or (layer0_outputs(1020)));
    outputs(495) <= not(layer0_outputs(856));
    outputs(496) <= '0';
    outputs(497) <= not((layer0_outputs(1014)) xor (layer0_outputs(1160)));
    outputs(498) <= not(layer0_outputs(2244));
    outputs(499) <= (layer0_outputs(1567)) and not (layer0_outputs(2413));
    outputs(500) <= not(layer0_outputs(1695));
    outputs(501) <= not((layer0_outputs(1819)) or (layer0_outputs(404)));
    outputs(502) <= (layer0_outputs(2045)) and (layer0_outputs(2180));
    outputs(503) <= not((layer0_outputs(1583)) or (layer0_outputs(491)));
    outputs(504) <= '0';
    outputs(505) <= layer0_outputs(1840);
    outputs(506) <= (layer0_outputs(1040)) and (layer0_outputs(610));
    outputs(507) <= not(layer0_outputs(347));
    outputs(508) <= layer0_outputs(1157);
    outputs(509) <= not((layer0_outputs(1095)) xor (layer0_outputs(227)));
    outputs(510) <= (layer0_outputs(1068)) and not (layer0_outputs(2398));
    outputs(511) <= not(layer0_outputs(180));
    outputs(512) <= layer0_outputs(2172);
    outputs(513) <= (layer0_outputs(1277)) xor (layer0_outputs(624));
    outputs(514) <= layer0_outputs(1121);
    outputs(515) <= not((layer0_outputs(763)) or (layer0_outputs(2541)));
    outputs(516) <= not(layer0_outputs(737));
    outputs(517) <= not((layer0_outputs(626)) or (layer0_outputs(1226)));
    outputs(518) <= layer0_outputs(2325);
    outputs(519) <= not((layer0_outputs(245)) xor (layer0_outputs(1351)));
    outputs(520) <= not((layer0_outputs(1891)) xor (layer0_outputs(206)));
    outputs(521) <= layer0_outputs(2522);
    outputs(522) <= not(layer0_outputs(947));
    outputs(523) <= not(layer0_outputs(2014));
    outputs(524) <= layer0_outputs(2314);
    outputs(525) <= layer0_outputs(1401);
    outputs(526) <= (layer0_outputs(2250)) and not (layer0_outputs(777));
    outputs(527) <= not(layer0_outputs(341));
    outputs(528) <= (layer0_outputs(850)) and not (layer0_outputs(1646));
    outputs(529) <= not(layer0_outputs(1771));
    outputs(530) <= not(layer0_outputs(2030));
    outputs(531) <= layer0_outputs(1575);
    outputs(532) <= layer0_outputs(82);
    outputs(533) <= layer0_outputs(128);
    outputs(534) <= not((layer0_outputs(229)) xor (layer0_outputs(1935)));
    outputs(535) <= not(layer0_outputs(1945));
    outputs(536) <= not(layer0_outputs(2261)) or (layer0_outputs(2558));
    outputs(537) <= not(layer0_outputs(909)) or (layer0_outputs(1725));
    outputs(538) <= not(layer0_outputs(362));
    outputs(539) <= not(layer0_outputs(1902));
    outputs(540) <= not(layer0_outputs(424));
    outputs(541) <= not(layer0_outputs(1752));
    outputs(542) <= not((layer0_outputs(2457)) xor (layer0_outputs(415)));
    outputs(543) <= layer0_outputs(2242);
    outputs(544) <= (layer0_outputs(59)) xor (layer0_outputs(658));
    outputs(545) <= layer0_outputs(1482);
    outputs(546) <= layer0_outputs(2109);
    outputs(547) <= not(layer0_outputs(542)) or (layer0_outputs(1927));
    outputs(548) <= not(layer0_outputs(656)) or (layer0_outputs(254));
    outputs(549) <= layer0_outputs(337);
    outputs(550) <= not(layer0_outputs(36)) or (layer0_outputs(1249));
    outputs(551) <= (layer0_outputs(132)) or (layer0_outputs(1378));
    outputs(552) <= layer0_outputs(1082);
    outputs(553) <= '1';
    outputs(554) <= not((layer0_outputs(579)) and (layer0_outputs(2107)));
    outputs(555) <= (layer0_outputs(1542)) and not (layer0_outputs(459));
    outputs(556) <= (layer0_outputs(1246)) or (layer0_outputs(2474));
    outputs(557) <= layer0_outputs(2546);
    outputs(558) <= not((layer0_outputs(442)) or (layer0_outputs(719)));
    outputs(559) <= not((layer0_outputs(355)) and (layer0_outputs(1046)));
    outputs(560) <= not((layer0_outputs(1878)) and (layer0_outputs(1770)));
    outputs(561) <= (layer0_outputs(1620)) xor (layer0_outputs(2468));
    outputs(562) <= not(layer0_outputs(1018));
    outputs(563) <= not(layer0_outputs(2530)) or (layer0_outputs(384));
    outputs(564) <= layer0_outputs(1340);
    outputs(565) <= layer0_outputs(476);
    outputs(566) <= layer0_outputs(350);
    outputs(567) <= not(layer0_outputs(1216));
    outputs(568) <= layer0_outputs(1521);
    outputs(569) <= not(layer0_outputs(2128));
    outputs(570) <= not(layer0_outputs(65));
    outputs(571) <= (layer0_outputs(2109)) and (layer0_outputs(2523));
    outputs(572) <= not(layer0_outputs(1197)) or (layer0_outputs(489));
    outputs(573) <= (layer0_outputs(1067)) xor (layer0_outputs(2065));
    outputs(574) <= layer0_outputs(1487);
    outputs(575) <= layer0_outputs(686);
    outputs(576) <= (layer0_outputs(2197)) or (layer0_outputs(1440));
    outputs(577) <= layer0_outputs(1703);
    outputs(578) <= layer0_outputs(401);
    outputs(579) <= not((layer0_outputs(2127)) and (layer0_outputs(1693)));
    outputs(580) <= layer0_outputs(212);
    outputs(581) <= layer0_outputs(525);
    outputs(582) <= not((layer0_outputs(1235)) or (layer0_outputs(487)));
    outputs(583) <= not(layer0_outputs(567));
    outputs(584) <= '1';
    outputs(585) <= (layer0_outputs(491)) xor (layer0_outputs(2375));
    outputs(586) <= not((layer0_outputs(1854)) or (layer0_outputs(1921)));
    outputs(587) <= layer0_outputs(1468);
    outputs(588) <= (layer0_outputs(1943)) and not (layer0_outputs(1536));
    outputs(589) <= layer0_outputs(2214);
    outputs(590) <= not((layer0_outputs(903)) or (layer0_outputs(2436)));
    outputs(591) <= not(layer0_outputs(726)) or (layer0_outputs(1374));
    outputs(592) <= layer0_outputs(899);
    outputs(593) <= not(layer0_outputs(219));
    outputs(594) <= (layer0_outputs(467)) and not (layer0_outputs(1411));
    outputs(595) <= (layer0_outputs(452)) or (layer0_outputs(425));
    outputs(596) <= not(layer0_outputs(1506));
    outputs(597) <= not((layer0_outputs(1662)) or (layer0_outputs(411)));
    outputs(598) <= not((layer0_outputs(58)) and (layer0_outputs(2031)));
    outputs(599) <= layer0_outputs(1323);
    outputs(600) <= not(layer0_outputs(535)) or (layer0_outputs(673));
    outputs(601) <= not(layer0_outputs(302)) or (layer0_outputs(1847));
    outputs(602) <= not(layer0_outputs(1949));
    outputs(603) <= not(layer0_outputs(135));
    outputs(604) <= not((layer0_outputs(444)) xor (layer0_outputs(685)));
    outputs(605) <= layer0_outputs(1406);
    outputs(606) <= not(layer0_outputs(1102));
    outputs(607) <= (layer0_outputs(2372)) and (layer0_outputs(1719));
    outputs(608) <= (layer0_outputs(756)) xor (layer0_outputs(2407));
    outputs(609) <= not(layer0_outputs(2487));
    outputs(610) <= not(layer0_outputs(1684)) or (layer0_outputs(244));
    outputs(611) <= not(layer0_outputs(1497));
    outputs(612) <= not((layer0_outputs(770)) and (layer0_outputs(201)));
    outputs(613) <= layer0_outputs(326);
    outputs(614) <= (layer0_outputs(2066)) xor (layer0_outputs(1648));
    outputs(615) <= not(layer0_outputs(728));
    outputs(616) <= (layer0_outputs(868)) and not (layer0_outputs(1415));
    outputs(617) <= not((layer0_outputs(339)) xor (layer0_outputs(2048)));
    outputs(618) <= not(layer0_outputs(2465));
    outputs(619) <= layer0_outputs(1954);
    outputs(620) <= not(layer0_outputs(71));
    outputs(621) <= (layer0_outputs(357)) or (layer0_outputs(458));
    outputs(622) <= not(layer0_outputs(2156));
    outputs(623) <= (layer0_outputs(1152)) and not (layer0_outputs(80));
    outputs(624) <= layer0_outputs(1049);
    outputs(625) <= (layer0_outputs(472)) or (layer0_outputs(2286));
    outputs(626) <= not((layer0_outputs(16)) or (layer0_outputs(1888)));
    outputs(627) <= not((layer0_outputs(2202)) and (layer0_outputs(1361)));
    outputs(628) <= not(layer0_outputs(195));
    outputs(629) <= (layer0_outputs(1593)) and (layer0_outputs(2372));
    outputs(630) <= (layer0_outputs(1091)) xor (layer0_outputs(996));
    outputs(631) <= not((layer0_outputs(2164)) and (layer0_outputs(2116)));
    outputs(632) <= not(layer0_outputs(2481));
    outputs(633) <= (layer0_outputs(1355)) and not (layer0_outputs(2450));
    outputs(634) <= not(layer0_outputs(1675)) or (layer0_outputs(1565));
    outputs(635) <= not((layer0_outputs(1566)) or (layer0_outputs(633)));
    outputs(636) <= (layer0_outputs(524)) xor (layer0_outputs(1063));
    outputs(637) <= not((layer0_outputs(1834)) and (layer0_outputs(1075)));
    outputs(638) <= not(layer0_outputs(2058));
    outputs(639) <= not((layer0_outputs(96)) and (layer0_outputs(587)));
    outputs(640) <= not((layer0_outputs(2323)) xor (layer0_outputs(2026)));
    outputs(641) <= layer0_outputs(1244);
    outputs(642) <= not((layer0_outputs(241)) or (layer0_outputs(192)));
    outputs(643) <= layer0_outputs(1876);
    outputs(644) <= not(layer0_outputs(1048));
    outputs(645) <= layer0_outputs(1918);
    outputs(646) <= (layer0_outputs(821)) xor (layer0_outputs(1726));
    outputs(647) <= (layer0_outputs(1100)) xor (layer0_outputs(1008));
    outputs(648) <= not(layer0_outputs(1435));
    outputs(649) <= not((layer0_outputs(2557)) or (layer0_outputs(2526)));
    outputs(650) <= not((layer0_outputs(1478)) or (layer0_outputs(1024)));
    outputs(651) <= layer0_outputs(2535);
    outputs(652) <= not(layer0_outputs(2543));
    outputs(653) <= not((layer0_outputs(1576)) and (layer0_outputs(2185)));
    outputs(654) <= not((layer0_outputs(1059)) and (layer0_outputs(1156)));
    outputs(655) <= not((layer0_outputs(1293)) and (layer0_outputs(838)));
    outputs(656) <= not((layer0_outputs(977)) xor (layer0_outputs(2215)));
    outputs(657) <= not((layer0_outputs(1278)) xor (layer0_outputs(1861)));
    outputs(658) <= layer0_outputs(607);
    outputs(659) <= not((layer0_outputs(1774)) or (layer0_outputs(464)));
    outputs(660) <= not(layer0_outputs(2009)) or (layer0_outputs(1860));
    outputs(661) <= (layer0_outputs(2280)) xor (layer0_outputs(296));
    outputs(662) <= not((layer0_outputs(154)) xor (layer0_outputs(173)));
    outputs(663) <= not(layer0_outputs(202)) or (layer0_outputs(1301));
    outputs(664) <= not(layer0_outputs(2102));
    outputs(665) <= not(layer0_outputs(555));
    outputs(666) <= not((layer0_outputs(85)) and (layer0_outputs(1835)));
    outputs(667) <= (layer0_outputs(1580)) or (layer0_outputs(1403));
    outputs(668) <= not(layer0_outputs(1754)) or (layer0_outputs(233));
    outputs(669) <= not(layer0_outputs(2349)) or (layer0_outputs(212));
    outputs(670) <= not((layer0_outputs(1232)) and (layer0_outputs(426)));
    outputs(671) <= layer0_outputs(2326);
    outputs(672) <= not((layer0_outputs(1533)) or (layer0_outputs(2154)));
    outputs(673) <= not(layer0_outputs(2410)) or (layer0_outputs(1594));
    outputs(674) <= not(layer0_outputs(2439)) or (layer0_outputs(1778));
    outputs(675) <= not(layer0_outputs(709));
    outputs(676) <= not((layer0_outputs(514)) and (layer0_outputs(2504)));
    outputs(677) <= (layer0_outputs(2000)) xor (layer0_outputs(1489));
    outputs(678) <= layer0_outputs(2063);
    outputs(679) <= not(layer0_outputs(873));
    outputs(680) <= not((layer0_outputs(2427)) xor (layer0_outputs(343)));
    outputs(681) <= not(layer0_outputs(1089)) or (layer0_outputs(2344));
    outputs(682) <= not((layer0_outputs(215)) and (layer0_outputs(2163)));
    outputs(683) <= not(layer0_outputs(1901));
    outputs(684) <= layer0_outputs(1572);
    outputs(685) <= not(layer0_outputs(162));
    outputs(686) <= not(layer0_outputs(566)) or (layer0_outputs(1875));
    outputs(687) <= (layer0_outputs(1427)) or (layer0_outputs(2429));
    outputs(688) <= not((layer0_outputs(2506)) xor (layer0_outputs(1841)));
    outputs(689) <= not(layer0_outputs(1925));
    outputs(690) <= (layer0_outputs(1135)) xor (layer0_outputs(1500));
    outputs(691) <= (layer0_outputs(1816)) and not (layer0_outputs(2499));
    outputs(692) <= not(layer0_outputs(1271));
    outputs(693) <= (layer0_outputs(494)) and not (layer0_outputs(216));
    outputs(694) <= not(layer0_outputs(923)) or (layer0_outputs(1971));
    outputs(695) <= not(layer0_outputs(1250));
    outputs(696) <= layer0_outputs(2038);
    outputs(697) <= not((layer0_outputs(2434)) or (layer0_outputs(1774)));
    outputs(698) <= not(layer0_outputs(903)) or (layer0_outputs(2371));
    outputs(699) <= not(layer0_outputs(1552)) or (layer0_outputs(292));
    outputs(700) <= not(layer0_outputs(269));
    outputs(701) <= layer0_outputs(570);
    outputs(702) <= layer0_outputs(672);
    outputs(703) <= not((layer0_outputs(2194)) xor (layer0_outputs(447)));
    outputs(704) <= not(layer0_outputs(53));
    outputs(705) <= (layer0_outputs(2478)) and (layer0_outputs(800));
    outputs(706) <= not(layer0_outputs(140)) or (layer0_outputs(768));
    outputs(707) <= layer0_outputs(1993);
    outputs(708) <= not((layer0_outputs(538)) xor (layer0_outputs(2076)));
    outputs(709) <= (layer0_outputs(899)) or (layer0_outputs(792));
    outputs(710) <= layer0_outputs(2230);
    outputs(711) <= not((layer0_outputs(811)) xor (layer0_outputs(891)));
    outputs(712) <= (layer0_outputs(1053)) and not (layer0_outputs(1220));
    outputs(713) <= not((layer0_outputs(634)) and (layer0_outputs(2051)));
    outputs(714) <= not(layer0_outputs(1787));
    outputs(715) <= (layer0_outputs(1054)) or (layer0_outputs(1319));
    outputs(716) <= (layer0_outputs(812)) xor (layer0_outputs(97));
    outputs(717) <= layer0_outputs(2142);
    outputs(718) <= layer0_outputs(2132);
    outputs(719) <= (layer0_outputs(2352)) or (layer0_outputs(1709));
    outputs(720) <= not(layer0_outputs(995));
    outputs(721) <= layer0_outputs(1763);
    outputs(722) <= (layer0_outputs(1893)) and not (layer0_outputs(2275));
    outputs(723) <= layer0_outputs(669);
    outputs(724) <= not(layer0_outputs(639));
    outputs(725) <= not(layer0_outputs(370));
    outputs(726) <= not((layer0_outputs(2189)) and (layer0_outputs(1596)));
    outputs(727) <= not((layer0_outputs(1938)) and (layer0_outputs(2149)));
    outputs(728) <= not((layer0_outputs(57)) or (layer0_outputs(440)));
    outputs(729) <= (layer0_outputs(1422)) and not (layer0_outputs(1747));
    outputs(730) <= not(layer0_outputs(1835));
    outputs(731) <= not(layer0_outputs(2196));
    outputs(732) <= layer0_outputs(1083);
    outputs(733) <= layer0_outputs(864);
    outputs(734) <= (layer0_outputs(159)) or (layer0_outputs(393));
    outputs(735) <= not(layer0_outputs(47));
    outputs(736) <= not(layer0_outputs(1096)) or (layer0_outputs(2309));
    outputs(737) <= not(layer0_outputs(2160)) or (layer0_outputs(329));
    outputs(738) <= not(layer0_outputs(1212)) or (layer0_outputs(409));
    outputs(739) <= (layer0_outputs(1658)) and not (layer0_outputs(1797));
    outputs(740) <= not((layer0_outputs(620)) or (layer0_outputs(1827)));
    outputs(741) <= layer0_outputs(1103);
    outputs(742) <= not(layer0_outputs(1383)) or (layer0_outputs(999));
    outputs(743) <= not(layer0_outputs(592)) or (layer0_outputs(881));
    outputs(744) <= (layer0_outputs(1837)) or (layer0_outputs(2022));
    outputs(745) <= layer0_outputs(2475);
    outputs(746) <= not(layer0_outputs(549));
    outputs(747) <= not(layer0_outputs(514));
    outputs(748) <= not(layer0_outputs(10));
    outputs(749) <= not(layer0_outputs(1558));
    outputs(750) <= layer0_outputs(882);
    outputs(751) <= (layer0_outputs(1379)) or (layer0_outputs(149));
    outputs(752) <= layer0_outputs(799);
    outputs(753) <= (layer0_outputs(1469)) xor (layer0_outputs(2215));
    outputs(754) <= layer0_outputs(1318);
    outputs(755) <= layer0_outputs(1511);
    outputs(756) <= not((layer0_outputs(581)) or (layer0_outputs(1383)));
    outputs(757) <= not(layer0_outputs(1907));
    outputs(758) <= (layer0_outputs(1316)) xor (layer0_outputs(1097));
    outputs(759) <= not(layer0_outputs(1809));
    outputs(760) <= not(layer0_outputs(122));
    outputs(761) <= (layer0_outputs(334)) and not (layer0_outputs(2170));
    outputs(762) <= layer0_outputs(2054);
    outputs(763) <= (layer0_outputs(2553)) and (layer0_outputs(1626));
    outputs(764) <= (layer0_outputs(2228)) xor (layer0_outputs(101));
    outputs(765) <= not(layer0_outputs(1296));
    outputs(766) <= not(layer0_outputs(602));
    outputs(767) <= not(layer0_outputs(1781));
    outputs(768) <= (layer0_outputs(2509)) and not (layer0_outputs(1212));
    outputs(769) <= layer0_outputs(652);
    outputs(770) <= layer0_outputs(2424);
    outputs(771) <= (layer0_outputs(1443)) xor (layer0_outputs(1424));
    outputs(772) <= (layer0_outputs(1814)) xor (layer0_outputs(2297));
    outputs(773) <= not(layer0_outputs(111));
    outputs(774) <= (layer0_outputs(57)) and (layer0_outputs(1320));
    outputs(775) <= (layer0_outputs(710)) xor (layer0_outputs(1914));
    outputs(776) <= (layer0_outputs(2252)) or (layer0_outputs(528));
    outputs(777) <= layer0_outputs(86);
    outputs(778) <= not(layer0_outputs(1236));
    outputs(779) <= (layer0_outputs(1987)) and not (layer0_outputs(1999));
    outputs(780) <= (layer0_outputs(1995)) or (layer0_outputs(1762));
    outputs(781) <= not(layer0_outputs(145));
    outputs(782) <= not(layer0_outputs(553)) or (layer0_outputs(663));
    outputs(783) <= not((layer0_outputs(162)) or (layer0_outputs(1586)));
    outputs(784) <= layer0_outputs(2115);
    outputs(785) <= not(layer0_outputs(822)) or (layer0_outputs(1758));
    outputs(786) <= layer0_outputs(613);
    outputs(787) <= not(layer0_outputs(1808));
    outputs(788) <= (layer0_outputs(2278)) and not (layer0_outputs(1632));
    outputs(789) <= (layer0_outputs(1413)) xor (layer0_outputs(1431));
    outputs(790) <= not(layer0_outputs(236));
    outputs(791) <= layer0_outputs(928);
    outputs(792) <= layer0_outputs(1644);
    outputs(793) <= not((layer0_outputs(106)) xor (layer0_outputs(2446)));
    outputs(794) <= (layer0_outputs(684)) and not (layer0_outputs(55));
    outputs(795) <= not(layer0_outputs(1894)) or (layer0_outputs(906));
    outputs(796) <= (layer0_outputs(1880)) xor (layer0_outputs(1430));
    outputs(797) <= (layer0_outputs(680)) xor (layer0_outputs(1671));
    outputs(798) <= (layer0_outputs(1571)) xor (layer0_outputs(2206));
    outputs(799) <= not(layer0_outputs(1793));
    outputs(800) <= not(layer0_outputs(1335)) or (layer0_outputs(2358));
    outputs(801) <= (layer0_outputs(1483)) or (layer0_outputs(617));
    outputs(802) <= layer0_outputs(2024);
    outputs(803) <= not(layer0_outputs(404)) or (layer0_outputs(559));
    outputs(804) <= (layer0_outputs(1737)) or (layer0_outputs(2043));
    outputs(805) <= layer0_outputs(1084);
    outputs(806) <= not(layer0_outputs(1429));
    outputs(807) <= (layer0_outputs(1435)) xor (layer0_outputs(992));
    outputs(808) <= not(layer0_outputs(1506));
    outputs(809) <= not(layer0_outputs(1538));
    outputs(810) <= layer0_outputs(1363);
    outputs(811) <= not((layer0_outputs(2110)) or (layer0_outputs(1627)));
    outputs(812) <= not(layer0_outputs(1624));
    outputs(813) <= layer0_outputs(627);
    outputs(814) <= layer0_outputs(1591);
    outputs(815) <= (layer0_outputs(493)) and (layer0_outputs(2320));
    outputs(816) <= layer0_outputs(2209);
    outputs(817) <= not(layer0_outputs(313));
    outputs(818) <= not(layer0_outputs(2419));
    outputs(819) <= not(layer0_outputs(1848));
    outputs(820) <= (layer0_outputs(807)) xor (layer0_outputs(2042));
    outputs(821) <= not((layer0_outputs(5)) xor (layer0_outputs(1036)));
    outputs(822) <= not((layer0_outputs(416)) and (layer0_outputs(609)));
    outputs(823) <= (layer0_outputs(2145)) and (layer0_outputs(601));
    outputs(824) <= not(layer0_outputs(1387));
    outputs(825) <= (layer0_outputs(1114)) and not (layer0_outputs(1012));
    outputs(826) <= not((layer0_outputs(884)) xor (layer0_outputs(562)));
    outputs(827) <= layer0_outputs(1740);
    outputs(828) <= not(layer0_outputs(1018));
    outputs(829) <= (layer0_outputs(1561)) and (layer0_outputs(2083));
    outputs(830) <= layer0_outputs(216);
    outputs(831) <= not(layer0_outputs(1563));
    outputs(832) <= layer0_outputs(407);
    outputs(833) <= (layer0_outputs(2406)) or (layer0_outputs(128));
    outputs(834) <= not(layer0_outputs(1182));
    outputs(835) <= not(layer0_outputs(1410));
    outputs(836) <= layer0_outputs(927);
    outputs(837) <= (layer0_outputs(2292)) and not (layer0_outputs(367));
    outputs(838) <= (layer0_outputs(701)) or (layer0_outputs(454));
    outputs(839) <= not(layer0_outputs(1642));
    outputs(840) <= (layer0_outputs(1396)) and (layer0_outputs(2114));
    outputs(841) <= (layer0_outputs(351)) or (layer0_outputs(674));
    outputs(842) <= (layer0_outputs(2032)) and (layer0_outputs(904));
    outputs(843) <= (layer0_outputs(1276)) and not (layer0_outputs(1180));
    outputs(844) <= layer0_outputs(1279);
    outputs(845) <= layer0_outputs(1655);
    outputs(846) <= layer0_outputs(681);
    outputs(847) <= not(layer0_outputs(648)) or (layer0_outputs(275));
    outputs(848) <= (layer0_outputs(787)) and not (layer0_outputs(2029));
    outputs(849) <= (layer0_outputs(1259)) and not (layer0_outputs(54));
    outputs(850) <= not(layer0_outputs(2313)) or (layer0_outputs(1398));
    outputs(851) <= (layer0_outputs(1077)) xor (layer0_outputs(564));
    outputs(852) <= (layer0_outputs(826)) or (layer0_outputs(2262));
    outputs(853) <= not((layer0_outputs(940)) and (layer0_outputs(997)));
    outputs(854) <= not((layer0_outputs(2165)) or (layer0_outputs(1910)));
    outputs(855) <= (layer0_outputs(1221)) or (layer0_outputs(1));
    outputs(856) <= not((layer0_outputs(2339)) or (layer0_outputs(1330)));
    outputs(857) <= not(layer0_outputs(1546));
    outputs(858) <= layer0_outputs(183);
    outputs(859) <= layer0_outputs(508);
    outputs(860) <= layer0_outputs(2143);
    outputs(861) <= (layer0_outputs(1720)) and not (layer0_outputs(235));
    outputs(862) <= not((layer0_outputs(1765)) or (layer0_outputs(1976)));
    outputs(863) <= layer0_outputs(1475);
    outputs(864) <= not((layer0_outputs(463)) xor (layer0_outputs(1941)));
    outputs(865) <= not(layer0_outputs(621));
    outputs(866) <= not(layer0_outputs(2153)) or (layer0_outputs(953));
    outputs(867) <= not((layer0_outputs(2345)) or (layer0_outputs(1734)));
    outputs(868) <= layer0_outputs(414);
    outputs(869) <= not(layer0_outputs(2503));
    outputs(870) <= layer0_outputs(1920);
    outputs(871) <= not(layer0_outputs(1956));
    outputs(872) <= not(layer0_outputs(2256));
    outputs(873) <= layer0_outputs(465);
    outputs(874) <= layer0_outputs(2549);
    outputs(875) <= (layer0_outputs(563)) and not (layer0_outputs(1667));
    outputs(876) <= not(layer0_outputs(1155));
    outputs(877) <= (layer0_outputs(1471)) xor (layer0_outputs(2123));
    outputs(878) <= layer0_outputs(456);
    outputs(879) <= (layer0_outputs(345)) and not (layer0_outputs(1560));
    outputs(880) <= not(layer0_outputs(2411)) or (layer0_outputs(1940));
    outputs(881) <= (layer0_outputs(941)) and not (layer0_outputs(1107));
    outputs(882) <= not((layer0_outputs(1638)) xor (layer0_outputs(125)));
    outputs(883) <= (layer0_outputs(661)) and not (layer0_outputs(100));
    outputs(884) <= not((layer0_outputs(405)) and (layer0_outputs(950)));
    outputs(885) <= layer0_outputs(432);
    outputs(886) <= not((layer0_outputs(2399)) or (layer0_outputs(1734)));
    outputs(887) <= not((layer0_outputs(526)) xor (layer0_outputs(450)));
    outputs(888) <= layer0_outputs(1074);
    outputs(889) <= layer0_outputs(2182);
    outputs(890) <= not(layer0_outputs(40));
    outputs(891) <= (layer0_outputs(1686)) and not (layer0_outputs(1002));
    outputs(892) <= (layer0_outputs(811)) or (layer0_outputs(201));
    outputs(893) <= (layer0_outputs(1133)) and (layer0_outputs(1381));
    outputs(894) <= layer0_outputs(197);
    outputs(895) <= not(layer0_outputs(1268)) or (layer0_outputs(1043));
    outputs(896) <= layer0_outputs(1165);
    outputs(897) <= not(layer0_outputs(2173));
    outputs(898) <= not((layer0_outputs(1464)) xor (layer0_outputs(2521)));
    outputs(899) <= (layer0_outputs(2234)) xor (layer0_outputs(2158));
    outputs(900) <= not(layer0_outputs(1076));
    outputs(901) <= not(layer0_outputs(1229)) or (layer0_outputs(2479));
    outputs(902) <= not(layer0_outputs(548)) or (layer0_outputs(774));
    outputs(903) <= (layer0_outputs(531)) and not (layer0_outputs(306));
    outputs(904) <= not((layer0_outputs(263)) xor (layer0_outputs(2515)));
    outputs(905) <= (layer0_outputs(1951)) and (layer0_outputs(2177));
    outputs(906) <= not(layer0_outputs(920));
    outputs(907) <= not((layer0_outputs(2331)) and (layer0_outputs(469)));
    outputs(908) <= not(layer0_outputs(670));
    outputs(909) <= not((layer0_outputs(1604)) or (layer0_outputs(1491)));
    outputs(910) <= not((layer0_outputs(335)) xor (layer0_outputs(611)));
    outputs(911) <= layer0_outputs(2456);
    outputs(912) <= not(layer0_outputs(1231));
    outputs(913) <= not((layer0_outputs(843)) and (layer0_outputs(2253)));
    outputs(914) <= '1';
    outputs(915) <= not((layer0_outputs(322)) or (layer0_outputs(2233)));
    outputs(916) <= not((layer0_outputs(693)) xor (layer0_outputs(1977)));
    outputs(917) <= not(layer0_outputs(2401)) or (layer0_outputs(622));
    outputs(918) <= layer0_outputs(1074);
    outputs(919) <= (layer0_outputs(758)) and (layer0_outputs(214));
    outputs(920) <= not((layer0_outputs(379)) and (layer0_outputs(286)));
    outputs(921) <= (layer0_outputs(637)) xor (layer0_outputs(318));
    outputs(922) <= not((layer0_outputs(2064)) and (layer0_outputs(1973)));
    outputs(923) <= (layer0_outputs(660)) or (layer0_outputs(2118));
    outputs(924) <= layer0_outputs(939);
    outputs(925) <= not((layer0_outputs(2300)) or (layer0_outputs(1494)));
    outputs(926) <= (layer0_outputs(2166)) and not (layer0_outputs(116));
    outputs(927) <= not(layer0_outputs(930));
    outputs(928) <= not(layer0_outputs(1826));
    outputs(929) <= not(layer0_outputs(886));
    outputs(930) <= not((layer0_outputs(2357)) xor (layer0_outputs(153)));
    outputs(931) <= (layer0_outputs(917)) xor (layer0_outputs(727));
    outputs(932) <= (layer0_outputs(2431)) and (layer0_outputs(616));
    outputs(933) <= layer0_outputs(1281);
    outputs(934) <= not(layer0_outputs(1135)) or (layer0_outputs(1552));
    outputs(935) <= not(layer0_outputs(283));
    outputs(936) <= not((layer0_outputs(1796)) and (layer0_outputs(283)));
    outputs(937) <= (layer0_outputs(449)) xor (layer0_outputs(2285));
    outputs(938) <= (layer0_outputs(1276)) xor (layer0_outputs(1508));
    outputs(939) <= not(layer0_outputs(1391));
    outputs(940) <= layer0_outputs(2263);
    outputs(941) <= not((layer0_outputs(1125)) xor (layer0_outputs(67)));
    outputs(942) <= not((layer0_outputs(896)) xor (layer0_outputs(2379)));
    outputs(943) <= not((layer0_outputs(1401)) or (layer0_outputs(815)));
    outputs(944) <= not((layer0_outputs(2199)) or (layer0_outputs(1405)));
    outputs(945) <= not(layer0_outputs(184));
    outputs(946) <= not(layer0_outputs(914));
    outputs(947) <= not(layer0_outputs(236));
    outputs(948) <= (layer0_outputs(1441)) and (layer0_outputs(739));
    outputs(949) <= '1';
    outputs(950) <= not((layer0_outputs(2306)) xor (layer0_outputs(1993)));
    outputs(951) <= not((layer0_outputs(1584)) and (layer0_outputs(136)));
    outputs(952) <= (layer0_outputs(1908)) and not (layer0_outputs(88));
    outputs(953) <= not(layer0_outputs(1632));
    outputs(954) <= (layer0_outputs(2013)) or (layer0_outputs(1670));
    outputs(955) <= (layer0_outputs(2426)) and (layer0_outputs(1598));
    outputs(956) <= not((layer0_outputs(1479)) xor (layer0_outputs(1385)));
    outputs(957) <= layer0_outputs(1547);
    outputs(958) <= not(layer0_outputs(1913));
    outputs(959) <= not(layer0_outputs(2009)) or (layer0_outputs(2409));
    outputs(960) <= not(layer0_outputs(1392));
    outputs(961) <= not(layer0_outputs(1874)) or (layer0_outputs(2226));
    outputs(962) <= not(layer0_outputs(376));
    outputs(963) <= not(layer0_outputs(1206));
    outputs(964) <= (layer0_outputs(2182)) and not (layer0_outputs(894));
    outputs(965) <= (layer0_outputs(1336)) and not (layer0_outputs(2291));
    outputs(966) <= (layer0_outputs(1462)) or (layer0_outputs(2249));
    outputs(967) <= (layer0_outputs(2349)) xor (layer0_outputs(2148));
    outputs(968) <= (layer0_outputs(1660)) and not (layer0_outputs(848));
    outputs(969) <= layer0_outputs(716);
    outputs(970) <= (layer0_outputs(391)) and not (layer0_outputs(1205));
    outputs(971) <= (layer0_outputs(874)) or (layer0_outputs(862));
    outputs(972) <= not((layer0_outputs(1698)) or (layer0_outputs(40)));
    outputs(973) <= (layer0_outputs(157)) xor (layer0_outputs(172));
    outputs(974) <= (layer0_outputs(700)) or (layer0_outputs(2376));
    outputs(975) <= (layer0_outputs(113)) xor (layer0_outputs(2360));
    outputs(976) <= not((layer0_outputs(2292)) xor (layer0_outputs(1826)));
    outputs(977) <= not(layer0_outputs(1395));
    outputs(978) <= not(layer0_outputs(1351)) or (layer0_outputs(1839));
    outputs(979) <= not((layer0_outputs(78)) or (layer0_outputs(858)));
    outputs(980) <= not(layer0_outputs(977));
    outputs(981) <= not(layer0_outputs(1432));
    outputs(982) <= (layer0_outputs(1780)) and not (layer0_outputs(386));
    outputs(983) <= not((layer0_outputs(1969)) xor (layer0_outputs(950)));
    outputs(984) <= not(layer0_outputs(182));
    outputs(985) <= not((layer0_outputs(856)) or (layer0_outputs(948)));
    outputs(986) <= not((layer0_outputs(1579)) xor (layer0_outputs(609)));
    outputs(987) <= (layer0_outputs(2451)) and (layer0_outputs(1254));
    outputs(988) <= not(layer0_outputs(434));
    outputs(989) <= not(layer0_outputs(988)) or (layer0_outputs(2558));
    outputs(990) <= (layer0_outputs(1619)) or (layer0_outputs(2191));
    outputs(991) <= not((layer0_outputs(124)) and (layer0_outputs(1892)));
    outputs(992) <= not((layer0_outputs(859)) xor (layer0_outputs(931)));
    outputs(993) <= layer0_outputs(1313);
    outputs(994) <= layer0_outputs(28);
    outputs(995) <= (layer0_outputs(997)) and (layer0_outputs(546));
    outputs(996) <= layer0_outputs(1729);
    outputs(997) <= (layer0_outputs(1056)) and not (layer0_outputs(1880));
    outputs(998) <= (layer0_outputs(1958)) xor (layer0_outputs(2448));
    outputs(999) <= (layer0_outputs(1050)) or (layer0_outputs(1147));
    outputs(1000) <= layer0_outputs(1426);
    outputs(1001) <= (layer0_outputs(1312)) or (layer0_outputs(466));
    outputs(1002) <= (layer0_outputs(69)) xor (layer0_outputs(1428));
    outputs(1003) <= (layer0_outputs(223)) and not (layer0_outputs(2072));
    outputs(1004) <= layer0_outputs(1962);
    outputs(1005) <= layer0_outputs(265);
    outputs(1006) <= not((layer0_outputs(2021)) or (layer0_outputs(718)));
    outputs(1007) <= not(layer0_outputs(1712));
    outputs(1008) <= layer0_outputs(1763);
    outputs(1009) <= (layer0_outputs(1863)) or (layer0_outputs(678));
    outputs(1010) <= (layer0_outputs(696)) and not (layer0_outputs(101));
    outputs(1011) <= not(layer0_outputs(1356));
    outputs(1012) <= not((layer0_outputs(1003)) and (layer0_outputs(1623)));
    outputs(1013) <= layer0_outputs(1926);
    outputs(1014) <= (layer0_outputs(2356)) xor (layer0_outputs(18));
    outputs(1015) <= layer0_outputs(2159);
    outputs(1016) <= layer0_outputs(910);
    outputs(1017) <= not((layer0_outputs(1409)) or (layer0_outputs(121)));
    outputs(1018) <= not(layer0_outputs(620));
    outputs(1019) <= (layer0_outputs(985)) and (layer0_outputs(1818));
    outputs(1020) <= layer0_outputs(965);
    outputs(1021) <= layer0_outputs(2106);
    outputs(1022) <= not((layer0_outputs(671)) or (layer0_outputs(1438)));
    outputs(1023) <= (layer0_outputs(355)) or (layer0_outputs(2319));
    outputs(1024) <= layer0_outputs(665);
    outputs(1025) <= not((layer0_outputs(306)) xor (layer0_outputs(2061)));
    outputs(1026) <= not((layer0_outputs(2141)) and (layer0_outputs(60)));
    outputs(1027) <= (layer0_outputs(2519)) and not (layer0_outputs(393));
    outputs(1028) <= (layer0_outputs(2258)) xor (layer0_outputs(2235));
    outputs(1029) <= (layer0_outputs(905)) and not (layer0_outputs(2449));
    outputs(1030) <= (layer0_outputs(2380)) and not (layer0_outputs(1940));
    outputs(1031) <= not(layer0_outputs(276)) or (layer0_outputs(198));
    outputs(1032) <= (layer0_outputs(640)) and not (layer0_outputs(1407));
    outputs(1033) <= not(layer0_outputs(1694));
    outputs(1034) <= not((layer0_outputs(429)) or (layer0_outputs(2201)));
    outputs(1035) <= (layer0_outputs(73)) and not (layer0_outputs(1956));
    outputs(1036) <= not(layer0_outputs(560));
    outputs(1037) <= not(layer0_outputs(1355));
    outputs(1038) <= not(layer0_outputs(1731));
    outputs(1039) <= '0';
    outputs(1040) <= (layer0_outputs(323)) and not (layer0_outputs(1105));
    outputs(1041) <= (layer0_outputs(1828)) and (layer0_outputs(1369));
    outputs(1042) <= not(layer0_outputs(1947));
    outputs(1043) <= not((layer0_outputs(1917)) or (layer0_outputs(2444)));
    outputs(1044) <= (layer0_outputs(798)) and not (layer0_outputs(589));
    outputs(1045) <= (layer0_outputs(2531)) and (layer0_outputs(2282));
    outputs(1046) <= (layer0_outputs(765)) and not (layer0_outputs(1415));
    outputs(1047) <= not(layer0_outputs(2195));
    outputs(1048) <= not((layer0_outputs(1963)) or (layer0_outputs(645)));
    outputs(1049) <= (layer0_outputs(1333)) xor (layer0_outputs(684));
    outputs(1050) <= layer0_outputs(653);
    outputs(1051) <= not(layer0_outputs(1749));
    outputs(1052) <= (layer0_outputs(796)) and not (layer0_outputs(103));
    outputs(1053) <= not(layer0_outputs(1856));
    outputs(1054) <= not((layer0_outputs(734)) or (layer0_outputs(1899)));
    outputs(1055) <= (layer0_outputs(969)) and not (layer0_outputs(1330));
    outputs(1056) <= not(layer0_outputs(699));
    outputs(1057) <= (layer0_outputs(1146)) and (layer0_outputs(185));
    outputs(1058) <= (layer0_outputs(1166)) and (layer0_outputs(1449));
    outputs(1059) <= layer0_outputs(1711);
    outputs(1060) <= layer0_outputs(446);
    outputs(1061) <= not(layer0_outputs(1821));
    outputs(1062) <= not((layer0_outputs(1329)) or (layer0_outputs(2145)));
    outputs(1063) <= (layer0_outputs(304)) and not (layer0_outputs(551));
    outputs(1064) <= not(layer0_outputs(1129));
    outputs(1065) <= (layer0_outputs(7)) xor (layer0_outputs(2540));
    outputs(1066) <= (layer0_outputs(613)) and not (layer0_outputs(2134));
    outputs(1067) <= (layer0_outputs(2540)) and not (layer0_outputs(1180));
    outputs(1068) <= not(layer0_outputs(791));
    outputs(1069) <= (layer0_outputs(1241)) and not (layer0_outputs(835));
    outputs(1070) <= not((layer0_outputs(248)) or (layer0_outputs(436)));
    outputs(1071) <= (layer0_outputs(1433)) and (layer0_outputs(2086));
    outputs(1072) <= (layer0_outputs(2018)) and not (layer0_outputs(628));
    outputs(1073) <= layer0_outputs(155);
    outputs(1074) <= layer0_outputs(930);
    outputs(1075) <= not((layer0_outputs(1194)) or (layer0_outputs(2496)));
    outputs(1076) <= layer0_outputs(880);
    outputs(1077) <= layer0_outputs(1376);
    outputs(1078) <= (layer0_outputs(1350)) or (layer0_outputs(529));
    outputs(1079) <= layer0_outputs(1512);
    outputs(1080) <= not(layer0_outputs(223)) or (layer0_outputs(835));
    outputs(1081) <= layer0_outputs(2389);
    outputs(1082) <= (layer0_outputs(1991)) and (layer0_outputs(1108));
    outputs(1083) <= (layer0_outputs(1913)) or (layer0_outputs(1578));
    outputs(1084) <= (layer0_outputs(1958)) and (layer0_outputs(2216));
    outputs(1085) <= layer0_outputs(2255);
    outputs(1086) <= (layer0_outputs(309)) and not (layer0_outputs(1033));
    outputs(1087) <= not(layer0_outputs(1196));
    outputs(1088) <= layer0_outputs(580);
    outputs(1089) <= (layer0_outputs(1713)) and not (layer0_outputs(918));
    outputs(1090) <= (layer0_outputs(1101)) and not (layer0_outputs(188));
    outputs(1091) <= not(layer0_outputs(1695));
    outputs(1092) <= layer0_outputs(194);
    outputs(1093) <= (layer0_outputs(29)) and (layer0_outputs(1872));
    outputs(1094) <= (layer0_outputs(949)) and not (layer0_outputs(682));
    outputs(1095) <= layer0_outputs(1983);
    outputs(1096) <= not((layer0_outputs(9)) and (layer0_outputs(2534)));
    outputs(1097) <= not(layer0_outputs(1272));
    outputs(1098) <= (layer0_outputs(687)) xor (layer0_outputs(1032));
    outputs(1099) <= not((layer0_outputs(1294)) xor (layer0_outputs(2467)));
    outputs(1100) <= (layer0_outputs(43)) and not (layer0_outputs(2151));
    outputs(1101) <= not((layer0_outputs(238)) or (layer0_outputs(644)));
    outputs(1102) <= (layer0_outputs(224)) and not (layer0_outputs(209));
    outputs(1103) <= not(layer0_outputs(1521)) or (layer0_outputs(1298));
    outputs(1104) <= (layer0_outputs(1051)) and not (layer0_outputs(21));
    outputs(1105) <= not((layer0_outputs(2121)) or (layer0_outputs(965)));
    outputs(1106) <= layer0_outputs(2186);
    outputs(1107) <= not((layer0_outputs(2425)) or (layer0_outputs(2220)));
    outputs(1108) <= layer0_outputs(580);
    outputs(1109) <= not((layer0_outputs(1178)) xor (layer0_outputs(957)));
    outputs(1110) <= (layer0_outputs(512)) and not (layer0_outputs(440));
    outputs(1111) <= (layer0_outputs(1626)) and (layer0_outputs(2173));
    outputs(1112) <= not(layer0_outputs(305));
    outputs(1113) <= layer0_outputs(737);
    outputs(1114) <= (layer0_outputs(2269)) and (layer0_outputs(1732));
    outputs(1115) <= layer0_outputs(1984);
    outputs(1116) <= (layer0_outputs(752)) and not (layer0_outputs(1243));
    outputs(1117) <= (layer0_outputs(741)) and (layer0_outputs(1314));
    outputs(1118) <= (layer0_outputs(2556)) and not (layer0_outputs(2362));
    outputs(1119) <= layer0_outputs(2021);
    outputs(1120) <= not((layer0_outputs(508)) or (layer0_outputs(1126)));
    outputs(1121) <= layer0_outputs(805);
    outputs(1122) <= not(layer0_outputs(1455));
    outputs(1123) <= layer0_outputs(502);
    outputs(1124) <= (layer0_outputs(1314)) and not (layer0_outputs(426));
    outputs(1125) <= not(layer0_outputs(455)) or (layer0_outputs(2204));
    outputs(1126) <= (layer0_outputs(439)) and not (layer0_outputs(1950));
    outputs(1127) <= not(layer0_outputs(74));
    outputs(1128) <= (layer0_outputs(22)) and not (layer0_outputs(1249));
    outputs(1129) <= not(layer0_outputs(328));
    outputs(1130) <= not(layer0_outputs(1300));
    outputs(1131) <= (layer0_outputs(304)) and not (layer0_outputs(831));
    outputs(1132) <= (layer0_outputs(1505)) and not (layer0_outputs(2124));
    outputs(1133) <= not(layer0_outputs(2547));
    outputs(1134) <= not(layer0_outputs(389));
    outputs(1135) <= not(layer0_outputs(525));
    outputs(1136) <= (layer0_outputs(1704)) or (layer0_outputs(1072));
    outputs(1137) <= (layer0_outputs(373)) and (layer0_outputs(1305));
    outputs(1138) <= layer0_outputs(916);
    outputs(1139) <= not(layer0_outputs(1636)) or (layer0_outputs(1198));
    outputs(1140) <= (layer0_outputs(1270)) and not (layer0_outputs(2329));
    outputs(1141) <= not(layer0_outputs(2350));
    outputs(1142) <= (layer0_outputs(2015)) and not (layer0_outputs(795));
    outputs(1143) <= (layer0_outputs(270)) and not (layer0_outputs(956));
    outputs(1144) <= not((layer0_outputs(482)) or (layer0_outputs(1654)));
    outputs(1145) <= layer0_outputs(239);
    outputs(1146) <= (layer0_outputs(629)) xor (layer0_outputs(976));
    outputs(1147) <= (layer0_outputs(1745)) and (layer0_outputs(1418));
    outputs(1148) <= layer0_outputs(221);
    outputs(1149) <= (layer0_outputs(1832)) and not (layer0_outputs(133));
    outputs(1150) <= not((layer0_outputs(1132)) or (layer0_outputs(1134)));
    outputs(1151) <= not(layer0_outputs(234)) or (layer0_outputs(1161));
    outputs(1152) <= not((layer0_outputs(586)) and (layer0_outputs(1058)));
    outputs(1153) <= (layer0_outputs(866)) xor (layer0_outputs(1796));
    outputs(1154) <= not(layer0_outputs(1290));
    outputs(1155) <= layer0_outputs(744);
    outputs(1156) <= (layer0_outputs(1005)) and not (layer0_outputs(933));
    outputs(1157) <= not((layer0_outputs(662)) xor (layer0_outputs(929)));
    outputs(1158) <= not((layer0_outputs(2329)) xor (layer0_outputs(138)));
    outputs(1159) <= not(layer0_outputs(1618));
    outputs(1160) <= layer0_outputs(853);
    outputs(1161) <= not(layer0_outputs(1265));
    outputs(1162) <= not((layer0_outputs(1918)) xor (layer0_outputs(708)));
    outputs(1163) <= (layer0_outputs(175)) and not (layer0_outputs(1564));
    outputs(1164) <= (layer0_outputs(2006)) and (layer0_outputs(246));
    outputs(1165) <= not((layer0_outputs(1017)) and (layer0_outputs(2236)));
    outputs(1166) <= not((layer0_outputs(574)) or (layer0_outputs(844)));
    outputs(1167) <= not(layer0_outputs(33));
    outputs(1168) <= not((layer0_outputs(2177)) xor (layer0_outputs(1924)));
    outputs(1169) <= (layer0_outputs(1054)) or (layer0_outputs(780));
    outputs(1170) <= not(layer0_outputs(2143));
    outputs(1171) <= (layer0_outputs(1325)) and not (layer0_outputs(158));
    outputs(1172) <= not(layer0_outputs(1683));
    outputs(1173) <= (layer0_outputs(97)) and (layer0_outputs(2528));
    outputs(1174) <= layer0_outputs(538);
    outputs(1175) <= not((layer0_outputs(1851)) or (layer0_outputs(2461)));
    outputs(1176) <= not(layer0_outputs(1454));
    outputs(1177) <= not(layer0_outputs(118));
    outputs(1178) <= not(layer0_outputs(1028));
    outputs(1179) <= layer0_outputs(1906);
    outputs(1180) <= layer0_outputs(863);
    outputs(1181) <= layer0_outputs(776);
    outputs(1182) <= not(layer0_outputs(2290));
    outputs(1183) <= (layer0_outputs(406)) and (layer0_outputs(2393));
    outputs(1184) <= (layer0_outputs(991)) and not (layer0_outputs(668));
    outputs(1185) <= (layer0_outputs(877)) and (layer0_outputs(1871));
    outputs(1186) <= (layer0_outputs(2488)) and not (layer0_outputs(866));
    outputs(1187) <= (layer0_outputs(667)) and not (layer0_outputs(385));
    outputs(1188) <= (layer0_outputs(309)) and (layer0_outputs(1464));
    outputs(1189) <= (layer0_outputs(595)) xor (layer0_outputs(922));
    outputs(1190) <= not((layer0_outputs(1030)) xor (layer0_outputs(2206)));
    outputs(1191) <= not((layer0_outputs(1755)) xor (layer0_outputs(627)));
    outputs(1192) <= layer0_outputs(281);
    outputs(1193) <= not(layer0_outputs(1382));
    outputs(1194) <= not(layer0_outputs(1006));
    outputs(1195) <= not(layer0_outputs(1866));
    outputs(1196) <= not(layer0_outputs(141));
    outputs(1197) <= (layer0_outputs(181)) and not (layer0_outputs(1768));
    outputs(1198) <= not((layer0_outputs(1104)) xor (layer0_outputs(1246)));
    outputs(1199) <= not(layer0_outputs(2284));
    outputs(1200) <= not(layer0_outputs(1137)) or (layer0_outputs(983));
    outputs(1201) <= (layer0_outputs(2417)) xor (layer0_outputs(416));
    outputs(1202) <= not((layer0_outputs(2161)) xor (layer0_outputs(2005)));
    outputs(1203) <= (layer0_outputs(1109)) xor (layer0_outputs(551));
    outputs(1204) <= layer0_outputs(1875);
    outputs(1205) <= (layer0_outputs(1073)) and not (layer0_outputs(1420));
    outputs(1206) <= (layer0_outputs(474)) and not (layer0_outputs(1300));
    outputs(1207) <= layer0_outputs(1000);
    outputs(1208) <= not(layer0_outputs(1685));
    outputs(1209) <= not(layer0_outputs(6));
    outputs(1210) <= not((layer0_outputs(2010)) or (layer0_outputs(507)));
    outputs(1211) <= (layer0_outputs(1206)) and not (layer0_outputs(2304));
    outputs(1212) <= not((layer0_outputs(2004)) or (layer0_outputs(2140)));
    outputs(1213) <= layer0_outputs(2482);
    outputs(1214) <= not((layer0_outputs(1923)) or (layer0_outputs(114)));
    outputs(1215) <= (layer0_outputs(539)) xor (layer0_outputs(970));
    outputs(1216) <= (layer0_outputs(762)) and (layer0_outputs(750));
    outputs(1217) <= not(layer0_outputs(1481));
    outputs(1218) <= not(layer0_outputs(418));
    outputs(1219) <= not((layer0_outputs(1944)) or (layer0_outputs(152)));
    outputs(1220) <= layer0_outputs(980);
    outputs(1221) <= not(layer0_outputs(259));
    outputs(1222) <= (layer0_outputs(2458)) and not (layer0_outputs(971));
    outputs(1223) <= (layer0_outputs(1584)) and not (layer0_outputs(2105));
    outputs(1224) <= '0';
    outputs(1225) <= layer0_outputs(936);
    outputs(1226) <= not((layer0_outputs(2433)) xor (layer0_outputs(2025)));
    outputs(1227) <= not(layer0_outputs(2245));
    outputs(1228) <= not((layer0_outputs(714)) or (layer0_outputs(1954)));
    outputs(1229) <= not((layer0_outputs(1264)) and (layer0_outputs(1718)));
    outputs(1230) <= (layer0_outputs(2354)) and not (layer0_outputs(71));
    outputs(1231) <= layer0_outputs(1750);
    outputs(1232) <= not((layer0_outputs(1557)) or (layer0_outputs(1998)));
    outputs(1233) <= not(layer0_outputs(1379));
    outputs(1234) <= layer0_outputs(1713);
    outputs(1235) <= not(layer0_outputs(532));
    outputs(1236) <= layer0_outputs(1833);
    outputs(1237) <= layer0_outputs(735);
    outputs(1238) <= (layer0_outputs(2138)) and (layer0_outputs(168));
    outputs(1239) <= not((layer0_outputs(1050)) or (layer0_outputs(1484)));
    outputs(1240) <= layer0_outputs(1000);
    outputs(1241) <= layer0_outputs(2012);
    outputs(1242) <= not(layer0_outputs(1690));
    outputs(1243) <= layer0_outputs(1430);
    outputs(1244) <= (layer0_outputs(1728)) xor (layer0_outputs(1630));
    outputs(1245) <= not((layer0_outputs(1553)) or (layer0_outputs(2232)));
    outputs(1246) <= not((layer0_outputs(1031)) or (layer0_outputs(2386)));
    outputs(1247) <= (layer0_outputs(827)) and (layer0_outputs(817));
    outputs(1248) <= layer0_outputs(2500);
    outputs(1249) <= not(layer0_outputs(1412));
    outputs(1250) <= not(layer0_outputs(1210));
    outputs(1251) <= layer0_outputs(1003);
    outputs(1252) <= (layer0_outputs(2484)) and not (layer0_outputs(60));
    outputs(1253) <= (layer0_outputs(517)) and not (layer0_outputs(1271));
    outputs(1254) <= not(layer0_outputs(2381));
    outputs(1255) <= (layer0_outputs(1543)) xor (layer0_outputs(1176));
    outputs(1256) <= (layer0_outputs(479)) and (layer0_outputs(1480));
    outputs(1257) <= not(layer0_outputs(2401));
    outputs(1258) <= layer0_outputs(2015);
    outputs(1259) <= layer0_outputs(2219);
    outputs(1260) <= not(layer0_outputs(348));
    outputs(1261) <= (layer0_outputs(889)) and not (layer0_outputs(2404));
    outputs(1262) <= (layer0_outputs(1260)) and (layer0_outputs(1245));
    outputs(1263) <= (layer0_outputs(2045)) and not (layer0_outputs(1526));
    outputs(1264) <= (layer0_outputs(1677)) xor (layer0_outputs(1555));
    outputs(1265) <= not((layer0_outputs(986)) or (layer0_outputs(2187)));
    outputs(1266) <= layer0_outputs(1410);
    outputs(1267) <= not((layer0_outputs(1683)) or (layer0_outputs(816)));
    outputs(1268) <= (layer0_outputs(608)) and not (layer0_outputs(1890));
    outputs(1269) <= (layer0_outputs(1512)) and not (layer0_outputs(1885));
    outputs(1270) <= not((layer0_outputs(1845)) xor (layer0_outputs(1966)));
    outputs(1271) <= (layer0_outputs(172)) and not (layer0_outputs(2053));
    outputs(1272) <= not((layer0_outputs(1928)) or (layer0_outputs(1299)));
    outputs(1273) <= not(layer0_outputs(1706)) or (layer0_outputs(906));
    outputs(1274) <= (layer0_outputs(1986)) and not (layer0_outputs(1932));
    outputs(1275) <= not(layer0_outputs(2322));
    outputs(1276) <= (layer0_outputs(1316)) and not (layer0_outputs(1953));
    outputs(1277) <= not(layer0_outputs(1643));
    outputs(1278) <= not(layer0_outputs(1822));
    outputs(1279) <= layer0_outputs(36);
    outputs(1280) <= not(layer0_outputs(2353)) or (layer0_outputs(2126));
    outputs(1281) <= layer0_outputs(932);
    outputs(1282) <= not((layer0_outputs(431)) and (layer0_outputs(1354)));
    outputs(1283) <= not(layer0_outputs(884));
    outputs(1284) <= (layer0_outputs(972)) xor (layer0_outputs(579));
    outputs(1285) <= not((layer0_outputs(781)) xor (layer0_outputs(1862)));
    outputs(1286) <= not(layer0_outputs(993)) or (layer0_outputs(2436));
    outputs(1287) <= not((layer0_outputs(993)) and (layer0_outputs(1795)));
    outputs(1288) <= (layer0_outputs(844)) or (layer0_outputs(1672));
    outputs(1289) <= not(layer0_outputs(1517));
    outputs(1290) <= layer0_outputs(1945);
    outputs(1291) <= '1';
    outputs(1292) <= not((layer0_outputs(1900)) xor (layer0_outputs(1665)));
    outputs(1293) <= not(layer0_outputs(2070));
    outputs(1294) <= not((layer0_outputs(865)) xor (layer0_outputs(1684)));
    outputs(1295) <= not((layer0_outputs(1533)) xor (layer0_outputs(1548)));
    outputs(1296) <= not((layer0_outputs(1442)) and (layer0_outputs(853)));
    outputs(1297) <= not(layer0_outputs(2463));
    outputs(1298) <= (layer0_outputs(2512)) xor (layer0_outputs(180));
    outputs(1299) <= not(layer0_outputs(1106));
    outputs(1300) <= not(layer0_outputs(1961));
    outputs(1301) <= (layer0_outputs(376)) xor (layer0_outputs(231));
    outputs(1302) <= (layer0_outputs(1477)) and (layer0_outputs(787));
    outputs(1303) <= not(layer0_outputs(1697));
    outputs(1304) <= layer0_outputs(1855);
    outputs(1305) <= (layer0_outputs(1419)) xor (layer0_outputs(2208));
    outputs(1306) <= not((layer0_outputs(183)) or (layer0_outputs(1200)));
    outputs(1307) <= layer0_outputs(1978);
    outputs(1308) <= not(layer0_outputs(257));
    outputs(1309) <= not((layer0_outputs(1140)) xor (layer0_outputs(456)));
    outputs(1310) <= (layer0_outputs(1927)) and (layer0_outputs(1191));
    outputs(1311) <= layer0_outputs(1498);
    outputs(1312) <= not((layer0_outputs(1573)) xor (layer0_outputs(1445)));
    outputs(1313) <= not(layer0_outputs(149));
    outputs(1314) <= (layer0_outputs(2344)) xor (layer0_outputs(729));
    outputs(1315) <= (layer0_outputs(1844)) xor (layer0_outputs(1142));
    outputs(1316) <= not(layer0_outputs(2205));
    outputs(1317) <= (layer0_outputs(381)) and not (layer0_outputs(177));
    outputs(1318) <= not((layer0_outputs(916)) and (layer0_outputs(983)));
    outputs(1319) <= not(layer0_outputs(1337));
    outputs(1320) <= not(layer0_outputs(156)) or (layer0_outputs(395));
    outputs(1321) <= not((layer0_outputs(1145)) xor (layer0_outputs(41)));
    outputs(1322) <= (layer0_outputs(501)) xor (layer0_outputs(1080));
    outputs(1323) <= layer0_outputs(511);
    outputs(1324) <= layer0_outputs(2246);
    outputs(1325) <= not(layer0_outputs(1873)) or (layer0_outputs(764));
    outputs(1326) <= layer0_outputs(608);
    outputs(1327) <= not(layer0_outputs(1037));
    outputs(1328) <= (layer0_outputs(2217)) and not (layer0_outputs(249));
    outputs(1329) <= not((layer0_outputs(2305)) xor (layer0_outputs(7)));
    outputs(1330) <= (layer0_outputs(687)) xor (layer0_outputs(1884));
    outputs(1331) <= (layer0_outputs(1293)) and (layer0_outputs(58));
    outputs(1332) <= (layer0_outputs(1640)) xor (layer0_outputs(2123));
    outputs(1333) <= (layer0_outputs(328)) or (layer0_outputs(471));
    outputs(1334) <= (layer0_outputs(427)) xor (layer0_outputs(1877));
    outputs(1335) <= not(layer0_outputs(2102)) or (layer0_outputs(1496));
    outputs(1336) <= (layer0_outputs(2049)) xor (layer0_outputs(1404));
    outputs(1337) <= layer0_outputs(1258);
    outputs(1338) <= (layer0_outputs(597)) xor (layer0_outputs(166));
    outputs(1339) <= not(layer0_outputs(1242));
    outputs(1340) <= not((layer0_outputs(641)) xor (layer0_outputs(2226)));
    outputs(1341) <= layer0_outputs(773);
    outputs(1342) <= not(layer0_outputs(1102)) or (layer0_outputs(1384));
    outputs(1343) <= (layer0_outputs(1611)) xor (layer0_outputs(1286));
    outputs(1344) <= (layer0_outputs(2207)) or (layer0_outputs(537));
    outputs(1345) <= not((layer0_outputs(412)) or (layer0_outputs(720)));
    outputs(1346) <= not(layer0_outputs(2139));
    outputs(1347) <= (layer0_outputs(2212)) xor (layer0_outputs(340));
    outputs(1348) <= not(layer0_outputs(955));
    outputs(1349) <= not(layer0_outputs(988)) or (layer0_outputs(49));
    outputs(1350) <= (layer0_outputs(1540)) and not (layer0_outputs(119));
    outputs(1351) <= (layer0_outputs(1955)) and not (layer0_outputs(1917));
    outputs(1352) <= (layer0_outputs(1612)) and not (layer0_outputs(570));
    outputs(1353) <= not((layer0_outputs(1762)) or (layer0_outputs(1083)));
    outputs(1354) <= layer0_outputs(1306);
    outputs(1355) <= layer0_outputs(926);
    outputs(1356) <= (layer0_outputs(2125)) and not (layer0_outputs(413));
    outputs(1357) <= not(layer0_outputs(2314));
    outputs(1358) <= not(layer0_outputs(319));
    outputs(1359) <= (layer0_outputs(779)) and not (layer0_outputs(1261));
    outputs(1360) <= (layer0_outputs(606)) xor (layer0_outputs(2334));
    outputs(1361) <= not(layer0_outputs(1472));
    outputs(1362) <= layer0_outputs(1776);
    outputs(1363) <= not(layer0_outputs(2260)) or (layer0_outputs(1921));
    outputs(1364) <= (layer0_outputs(702)) xor (layer0_outputs(715));
    outputs(1365) <= (layer0_outputs(2086)) and not (layer0_outputs(1957));
    outputs(1366) <= not(layer0_outputs(1181)) or (layer0_outputs(2334));
    outputs(1367) <= not((layer0_outputs(807)) xor (layer0_outputs(1664)));
    outputs(1368) <= not((layer0_outputs(1641)) xor (layer0_outputs(1671)));
    outputs(1369) <= layer0_outputs(2425);
    outputs(1370) <= (layer0_outputs(929)) and not (layer0_outputs(1625));
    outputs(1371) <= (layer0_outputs(584)) and (layer0_outputs(778));
    outputs(1372) <= (layer0_outputs(1256)) xor (layer0_outputs(1087));
    outputs(1373) <= not((layer0_outputs(710)) or (layer0_outputs(2242)));
    outputs(1374) <= (layer0_outputs(1988)) xor (layer0_outputs(731));
    outputs(1375) <= (layer0_outputs(1234)) xor (layer0_outputs(1326));
    outputs(1376) <= not(layer0_outputs(1830));
    outputs(1377) <= layer0_outputs(1456);
    outputs(1378) <= not(layer0_outputs(803));
    outputs(1379) <= not((layer0_outputs(859)) and (layer0_outputs(1745)));
    outputs(1380) <= not((layer0_outputs(1502)) xor (layer0_outputs(1548)));
    outputs(1381) <= (layer0_outputs(208)) xor (layer0_outputs(1045));
    outputs(1382) <= not((layer0_outputs(2088)) xor (layer0_outputs(763)));
    outputs(1383) <= not(layer0_outputs(2505));
    outputs(1384) <= not(layer0_outputs(2093));
    outputs(1385) <= layer0_outputs(1494);
    outputs(1386) <= (layer0_outputs(49)) xor (layer0_outputs(569));
    outputs(1387) <= not(layer0_outputs(2205));
    outputs(1388) <= not(layer0_outputs(375));
    outputs(1389) <= (layer0_outputs(765)) and (layer0_outputs(2438));
    outputs(1390) <= layer0_outputs(2281);
    outputs(1391) <= not((layer0_outputs(2185)) xor (layer0_outputs(2062)));
    outputs(1392) <= not((layer0_outputs(2020)) xor (layer0_outputs(1229)));
    outputs(1393) <= not(layer0_outputs(1154)) or (layer0_outputs(374));
    outputs(1394) <= layer0_outputs(2278);
    outputs(1395) <= layer0_outputs(1227);
    outputs(1396) <= not((layer0_outputs(1032)) and (layer0_outputs(2041)));
    outputs(1397) <= (layer0_outputs(1100)) and not (layer0_outputs(2074));
    outputs(1398) <= not(layer0_outputs(2108));
    outputs(1399) <= layer0_outputs(63);
    outputs(1400) <= (layer0_outputs(898)) and (layer0_outputs(1994));
    outputs(1401) <= layer0_outputs(2537);
    outputs(1402) <= not((layer0_outputs(1741)) xor (layer0_outputs(246)));
    outputs(1403) <= not((layer0_outputs(1935)) xor (layer0_outputs(522)));
    outputs(1404) <= (layer0_outputs(326)) and not (layer0_outputs(545));
    outputs(1405) <= not((layer0_outputs(1803)) or (layer0_outputs(1782)));
    outputs(1406) <= not((layer0_outputs(1493)) or (layer0_outputs(1448)));
    outputs(1407) <= (layer0_outputs(1279)) xor (layer0_outputs(117));
    outputs(1408) <= not(layer0_outputs(210));
    outputs(1409) <= (layer0_outputs(902)) and (layer0_outputs(1922));
    outputs(1410) <= layer0_outputs(655);
    outputs(1411) <= (layer0_outputs(262)) xor (layer0_outputs(1544));
    outputs(1412) <= not(layer0_outputs(1722));
    outputs(1413) <= not(layer0_outputs(239));
    outputs(1414) <= layer0_outputs(572);
    outputs(1415) <= (layer0_outputs(1607)) and not (layer0_outputs(2496));
    outputs(1416) <= (layer0_outputs(908)) and (layer0_outputs(2147));
    outputs(1417) <= not((layer0_outputs(1459)) xor (layer0_outputs(1265)));
    outputs(1418) <= layer0_outputs(1395);
    outputs(1419) <= (layer0_outputs(2105)) and (layer0_outputs(2047));
    outputs(1420) <= not((layer0_outputs(2494)) and (layer0_outputs(2183)));
    outputs(1421) <= (layer0_outputs(668)) or (layer0_outputs(268));
    outputs(1422) <= layer0_outputs(497);
    outputs(1423) <= layer0_outputs(735);
    outputs(1424) <= not((layer0_outputs(592)) xor (layer0_outputs(617)));
    outputs(1425) <= not((layer0_outputs(2400)) or (layer0_outputs(2368)));
    outputs(1426) <= not(layer0_outputs(2477));
    outputs(1427) <= (layer0_outputs(1215)) xor (layer0_outputs(473));
    outputs(1428) <= (layer0_outputs(2543)) and (layer0_outputs(211));
    outputs(1429) <= not((layer0_outputs(269)) xor (layer0_outputs(428)));
    outputs(1430) <= (layer0_outputs(1901)) and (layer0_outputs(2308));
    outputs(1431) <= (layer0_outputs(540)) and (layer0_outputs(1043));
    outputs(1432) <= (layer0_outputs(226)) and not (layer0_outputs(2538));
    outputs(1433) <= not(layer0_outputs(885));
    outputs(1434) <= not((layer0_outputs(683)) xor (layer0_outputs(1226)));
    outputs(1435) <= (layer0_outputs(828)) and (layer0_outputs(2317));
    outputs(1436) <= (layer0_outputs(2310)) xor (layer0_outputs(875));
    outputs(1437) <= (layer0_outputs(2041)) xor (layer0_outputs(1646));
    outputs(1438) <= layer0_outputs(2481);
    outputs(1439) <= not((layer0_outputs(1048)) or (layer0_outputs(188)));
    outputs(1440) <= not((layer0_outputs(1630)) and (layer0_outputs(1445)));
    outputs(1441) <= layer0_outputs(1616);
    outputs(1442) <= layer0_outputs(2408);
    outputs(1443) <= (layer0_outputs(245)) and not (layer0_outputs(2493));
    outputs(1444) <= (layer0_outputs(1239)) or (layer0_outputs(1975));
    outputs(1445) <= not(layer0_outputs(651)) or (layer0_outputs(1352));
    outputs(1446) <= layer0_outputs(65);
    outputs(1447) <= not(layer0_outputs(1026));
    outputs(1448) <= not(layer0_outputs(634));
    outputs(1449) <= layer0_outputs(2361);
    outputs(1450) <= layer0_outputs(141);
    outputs(1451) <= (layer0_outputs(401)) and not (layer0_outputs(1092));
    outputs(1452) <= layer0_outputs(1710);
    outputs(1453) <= layer0_outputs(1690);
    outputs(1454) <= not(layer0_outputs(1915));
    outputs(1455) <= layer0_outputs(330);
    outputs(1456) <= not(layer0_outputs(759));
    outputs(1457) <= not((layer0_outputs(2424)) xor (layer0_outputs(728)));
    outputs(1458) <= layer0_outputs(407);
    outputs(1459) <= not((layer0_outputs(337)) or (layer0_outputs(1916)));
    outputs(1460) <= (layer0_outputs(623)) xor (layer0_outputs(2362));
    outputs(1461) <= (layer0_outputs(1120)) and (layer0_outputs(1619));
    outputs(1462) <= not((layer0_outputs(2285)) and (layer0_outputs(1324)));
    outputs(1463) <= layer0_outputs(2219);
    outputs(1464) <= (layer0_outputs(1887)) and not (layer0_outputs(25));
    outputs(1465) <= not(layer0_outputs(934));
    outputs(1466) <= (layer0_outputs(587)) xor (layer0_outputs(2237));
    outputs(1467) <= layer0_outputs(1260);
    outputs(1468) <= (layer0_outputs(645)) and not (layer0_outputs(1765));
    outputs(1469) <= layer0_outputs(438);
    outputs(1470) <= (layer0_outputs(1283)) and (layer0_outputs(1159));
    outputs(1471) <= not((layer0_outputs(2061)) xor (layer0_outputs(382)));
    outputs(1472) <= not((layer0_outputs(1898)) xor (layer0_outputs(396)));
    outputs(1473) <= not(layer0_outputs(92)) or (layer0_outputs(1744));
    outputs(1474) <= not(layer0_outputs(469));
    outputs(1475) <= (layer0_outputs(2181)) xor (layer0_outputs(633));
    outputs(1476) <= not(layer0_outputs(403));
    outputs(1477) <= (layer0_outputs(398)) xor (layer0_outputs(556));
    outputs(1478) <= layer0_outputs(540);
    outputs(1479) <= not((layer0_outputs(2472)) xor (layer0_outputs(649)));
    outputs(1480) <= (layer0_outputs(1612)) and (layer0_outputs(1657));
    outputs(1481) <= not((layer0_outputs(2522)) xor (layer0_outputs(2234)));
    outputs(1482) <= layer0_outputs(909);
    outputs(1483) <= not(layer0_outputs(305));
    outputs(1484) <= layer0_outputs(612);
    outputs(1485) <= layer0_outputs(1247);
    outputs(1486) <= not((layer0_outputs(605)) or (layer0_outputs(1211)));
    outputs(1487) <= not((layer0_outputs(79)) xor (layer0_outputs(1881)));
    outputs(1488) <= (layer0_outputs(760)) and not (layer0_outputs(900));
    outputs(1489) <= (layer0_outputs(1820)) xor (layer0_outputs(2231));
    outputs(1490) <= not((layer0_outputs(2445)) xor (layer0_outputs(876)));
    outputs(1491) <= (layer0_outputs(1912)) xor (layer0_outputs(2306));
    outputs(1492) <= not((layer0_outputs(2172)) xor (layer0_outputs(1639)));
    outputs(1493) <= (layer0_outputs(2033)) xor (layer0_outputs(1079));
    outputs(1494) <= layer0_outputs(2119);
    outputs(1495) <= layer0_outputs(493);
    outputs(1496) <= not((layer0_outputs(1098)) xor (layer0_outputs(1539)));
    outputs(1497) <= (layer0_outputs(348)) and not (layer0_outputs(496));
    outputs(1498) <= layer0_outputs(267);
    outputs(1499) <= not((layer0_outputs(275)) or (layer0_outputs(360)));
    outputs(1500) <= (layer0_outputs(2380)) and not (layer0_outputs(2018));
    outputs(1501) <= not(layer0_outputs(1639));
    outputs(1502) <= not(layer0_outputs(37));
    outputs(1503) <= not(layer0_outputs(1450));
    outputs(1504) <= layer0_outputs(1440);
    outputs(1505) <= (layer0_outputs(642)) xor (layer0_outputs(2324));
    outputs(1506) <= layer0_outputs(1669);
    outputs(1507) <= (layer0_outputs(1015)) xor (layer0_outputs(998));
    outputs(1508) <= not(layer0_outputs(1962));
    outputs(1509) <= not(layer0_outputs(959)) or (layer0_outputs(2200));
    outputs(1510) <= not((layer0_outputs(1389)) xor (layer0_outputs(465)));
    outputs(1511) <= not(layer0_outputs(2513));
    outputs(1512) <= layer0_outputs(821);
    outputs(1513) <= (layer0_outputs(251)) xor (layer0_outputs(664));
    outputs(1514) <= not((layer0_outputs(2056)) xor (layer0_outputs(2094)));
    outputs(1515) <= (layer0_outputs(740)) xor (layer0_outputs(1176));
    outputs(1516) <= not(layer0_outputs(1542)) or (layer0_outputs(1139));
    outputs(1517) <= (layer0_outputs(1979)) and (layer0_outputs(753));
    outputs(1518) <= not(layer0_outputs(1346));
    outputs(1519) <= layer0_outputs(1362);
    outputs(1520) <= (layer0_outputs(510)) and not (layer0_outputs(1093));
    outputs(1521) <= not(layer0_outputs(544)) or (layer0_outputs(344));
    outputs(1522) <= not(layer0_outputs(1333));
    outputs(1523) <= layer0_outputs(395);
    outputs(1524) <= not(layer0_outputs(133));
    outputs(1525) <= (layer0_outputs(317)) and (layer0_outputs(516));
    outputs(1526) <= not(layer0_outputs(1961));
    outputs(1527) <= (layer0_outputs(84)) xor (layer0_outputs(784));
    outputs(1528) <= (layer0_outputs(382)) and not (layer0_outputs(643));
    outputs(1529) <= not(layer0_outputs(1393));
    outputs(1530) <= not((layer0_outputs(861)) xor (layer0_outputs(1647)));
    outputs(1531) <= not(layer0_outputs(2315));
    outputs(1532) <= (layer0_outputs(1858)) xor (layer0_outputs(979));
    outputs(1533) <= (layer0_outputs(654)) and (layer0_outputs(927));
    outputs(1534) <= not(layer0_outputs(2133));
    outputs(1535) <= layer0_outputs(1403);
    outputs(1536) <= layer0_outputs(198);
    outputs(1537) <= not((layer0_outputs(2283)) or (layer0_outputs(2517)));
    outputs(1538) <= not(layer0_outputs(1583));
    outputs(1539) <= not(layer0_outputs(498));
    outputs(1540) <= not((layer0_outputs(1930)) xor (layer0_outputs(1546)));
    outputs(1541) <= not(layer0_outputs(2504)) or (layer0_outputs(1904));
    outputs(1542) <= not(layer0_outputs(1554));
    outputs(1543) <= (layer0_outputs(2196)) xor (layer0_outputs(2377));
    outputs(1544) <= not(layer0_outputs(1283));
    outputs(1545) <= (layer0_outputs(1138)) and not (layer0_outputs(1701));
    outputs(1546) <= (layer0_outputs(1803)) xor (layer0_outputs(576));
    outputs(1547) <= not(layer0_outputs(2040)) or (layer0_outputs(1715));
    outputs(1548) <= not((layer0_outputs(1366)) xor (layer0_outputs(2492)));
    outputs(1549) <= (layer0_outputs(1336)) and not (layer0_outputs(2384));
    outputs(1550) <= not((layer0_outputs(814)) and (layer0_outputs(758)));
    outputs(1551) <= not(layer0_outputs(1077)) or (layer0_outputs(2548));
    outputs(1552) <= not(layer0_outputs(1213));
    outputs(1553) <= (layer0_outputs(190)) and not (layer0_outputs(2318));
    outputs(1554) <= (layer0_outputs(1486)) xor (layer0_outputs(913));
    outputs(1555) <= not(layer0_outputs(1130));
    outputs(1556) <= not(layer0_outputs(2058));
    outputs(1557) <= not((layer0_outputs(2062)) xor (layer0_outputs(1647)));
    outputs(1558) <= not((layer0_outputs(1688)) or (layer0_outputs(1787)));
    outputs(1559) <= not(layer0_outputs(2243));
    outputs(1560) <= (layer0_outputs(1718)) and not (layer0_outputs(678));
    outputs(1561) <= (layer0_outputs(2150)) and (layer0_outputs(2373));
    outputs(1562) <= not(layer0_outputs(883)) or (layer0_outputs(1617));
    outputs(1563) <= (layer0_outputs(1741)) and (layer0_outputs(1284));
    outputs(1564) <= (layer0_outputs(1865)) and (layer0_outputs(1622));
    outputs(1565) <= not(layer0_outputs(560));
    outputs(1566) <= layer0_outputs(531);
    outputs(1567) <= (layer0_outputs(2264)) xor (layer0_outputs(2027));
    outputs(1568) <= not(layer0_outputs(2267));
    outputs(1569) <= (layer0_outputs(1746)) xor (layer0_outputs(50));
    outputs(1570) <= not(layer0_outputs(604));
    outputs(1571) <= layer0_outputs(1503);
    outputs(1572) <= not((layer0_outputs(793)) or (layer0_outputs(1359)));
    outputs(1573) <= layer0_outputs(2270);
    outputs(1574) <= layer0_outputs(221);
    outputs(1575) <= not(layer0_outputs(2179)) or (layer0_outputs(483));
    outputs(1576) <= layer0_outputs(26);
    outputs(1577) <= (layer0_outputs(1380)) xor (layer0_outputs(1773));
    outputs(1578) <= not(layer0_outputs(1499)) or (layer0_outputs(1373));
    outputs(1579) <= not(layer0_outputs(2441));
    outputs(1580) <= (layer0_outputs(69)) and not (layer0_outputs(614));
    outputs(1581) <= layer0_outputs(195);
    outputs(1582) <= not(layer0_outputs(2338));
    outputs(1583) <= layer0_outputs(987);
    outputs(1584) <= (layer0_outputs(46)) and not (layer0_outputs(331));
    outputs(1585) <= layer0_outputs(1010);
    outputs(1586) <= layer0_outputs(2382);
    outputs(1587) <= not((layer0_outputs(1871)) xor (layer0_outputs(951)));
    outputs(1588) <= (layer0_outputs(1129)) and not (layer0_outputs(566));
    outputs(1589) <= layer0_outputs(1589);
    outputs(1590) <= not((layer0_outputs(2395)) or (layer0_outputs(922)));
    outputs(1591) <= (layer0_outputs(2068)) and not (layer0_outputs(619));
    outputs(1592) <= not((layer0_outputs(833)) xor (layer0_outputs(2130)));
    outputs(1593) <= (layer0_outputs(1568)) and not (layer0_outputs(226));
    outputs(1594) <= (layer0_outputs(2321)) xor (layer0_outputs(1674));
    outputs(1595) <= (layer0_outputs(1942)) xor (layer0_outputs(2010));
    outputs(1596) <= (layer0_outputs(1427)) and not (layer0_outputs(790));
    outputs(1597) <= layer0_outputs(278);
    outputs(1598) <= not((layer0_outputs(943)) and (layer0_outputs(2032)));
    outputs(1599) <= layer0_outputs(958);
    outputs(1600) <= layer0_outputs(1692);
    outputs(1601) <= not((layer0_outputs(2200)) or (layer0_outputs(2304)));
    outputs(1602) <= layer0_outputs(2400);
    outputs(1603) <= not(layer0_outputs(1824));
    outputs(1604) <= (layer0_outputs(1572)) xor (layer0_outputs(1305));
    outputs(1605) <= not(layer0_outputs(1842)) or (layer0_outputs(2348));
    outputs(1606) <= not((layer0_outputs(1814)) or (layer0_outputs(2268)));
    outputs(1607) <= (layer0_outputs(1929)) or (layer0_outputs(1586));
    outputs(1608) <= not((layer0_outputs(2218)) or (layer0_outputs(908)));
    outputs(1609) <= not((layer0_outputs(593)) and (layer0_outputs(86)));
    outputs(1610) <= layer0_outputs(1421);
    outputs(1611) <= not((layer0_outputs(586)) xor (layer0_outputs(1296)));
    outputs(1612) <= not(layer0_outputs(967));
    outputs(1613) <= not(layer0_outputs(2162));
    outputs(1614) <= (layer0_outputs(1287)) and not (layer0_outputs(2369));
    outputs(1615) <= (layer0_outputs(2414)) and not (layer0_outputs(1727));
    outputs(1616) <= not(layer0_outputs(1324));
    outputs(1617) <= (layer0_outputs(732)) and not (layer0_outputs(238));
    outputs(1618) <= not((layer0_outputs(616)) or (layer0_outputs(322)));
    outputs(1619) <= not(layer0_outputs(1117));
    outputs(1620) <= (layer0_outputs(2221)) or (layer0_outputs(176));
    outputs(1621) <= (layer0_outputs(647)) and (layer0_outputs(1310));
    outputs(1622) <= (layer0_outputs(2056)) or (layer0_outputs(2080));
    outputs(1623) <= not(layer0_outputs(904)) or (layer0_outputs(2194));
    outputs(1624) <= not((layer0_outputs(2541)) or (layer0_outputs(1872)));
    outputs(1625) <= not(layer0_outputs(2503)) or (layer0_outputs(1964));
    outputs(1626) <= layer0_outputs(705);
    outputs(1627) <= (layer0_outputs(1209)) and not (layer0_outputs(274));
    outputs(1628) <= (layer0_outputs(178)) and not (layer0_outputs(1571));
    outputs(1629) <= not((layer0_outputs(1709)) or (layer0_outputs(1354)));
    outputs(1630) <= layer0_outputs(2003);
    outputs(1631) <= not((layer0_outputs(736)) xor (layer0_outputs(1315)));
    outputs(1632) <= (layer0_outputs(559)) xor (layer0_outputs(1122));
    outputs(1633) <= '1';
    outputs(1634) <= (layer0_outputs(952)) and not (layer0_outputs(2409));
    outputs(1635) <= not(layer0_outputs(1870)) or (layer0_outputs(273));
    outputs(1636) <= (layer0_outputs(1779)) and not (layer0_outputs(358));
    outputs(1637) <= not((layer0_outputs(1620)) or (layer0_outputs(1791)));
    outputs(1638) <= (layer0_outputs(280)) xor (layer0_outputs(619));
    outputs(1639) <= (layer0_outputs(409)) and not (layer0_outputs(1504));
    outputs(1640) <= (layer0_outputs(591)) xor (layer0_outputs(1609));
    outputs(1641) <= not(layer0_outputs(2101));
    outputs(1642) <= layer0_outputs(1343);
    outputs(1643) <= not((layer0_outputs(792)) or (layer0_outputs(2510)));
    outputs(1644) <= layer0_outputs(1893);
    outputs(1645) <= not(layer0_outputs(1616));
    outputs(1646) <= (layer0_outputs(1810)) and not (layer0_outputs(1829));
    outputs(1647) <= not((layer0_outputs(2193)) or (layer0_outputs(2293)));
    outputs(1648) <= not(layer0_outputs(963));
    outputs(1649) <= not(layer0_outputs(175));
    outputs(1650) <= layer0_outputs(702);
    outputs(1651) <= not(layer0_outputs(631));
    outputs(1652) <= not((layer0_outputs(2467)) or (layer0_outputs(788)));
    outputs(1653) <= not(layer0_outputs(706));
    outputs(1654) <= not(layer0_outputs(558));
    outputs(1655) <= not(layer0_outputs(1700)) or (layer0_outputs(1345));
    outputs(1656) <= (layer0_outputs(1943)) and (layer0_outputs(402));
    outputs(1657) <= (layer0_outputs(1118)) xor (layer0_outputs(1253));
    outputs(1658) <= not(layer0_outputs(1851));
    outputs(1659) <= not(layer0_outputs(80));
    outputs(1660) <= not((layer0_outputs(2469)) or (layer0_outputs(942)));
    outputs(1661) <= not(layer0_outputs(1631));
    outputs(1662) <= not(layer0_outputs(312));
    outputs(1663) <= (layer0_outputs(786)) xor (layer0_outputs(151));
    outputs(1664) <= (layer0_outputs(661)) and (layer0_outputs(2432));
    outputs(1665) <= not(layer0_outputs(2294)) or (layer0_outputs(292));
    outputs(1666) <= (layer0_outputs(1016)) or (layer0_outputs(822));
    outputs(1667) <= (layer0_outputs(50)) and not (layer0_outputs(1495));
    outputs(1668) <= not((layer0_outputs(864)) xor (layer0_outputs(408)));
    outputs(1669) <= not((layer0_outputs(311)) or (layer0_outputs(1960)));
    outputs(1670) <= (layer0_outputs(521)) xor (layer0_outputs(954));
    outputs(1671) <= (layer0_outputs(2307)) and not (layer0_outputs(777));
    outputs(1672) <= not((layer0_outputs(697)) or (layer0_outputs(1638)));
    outputs(1673) <= layer0_outputs(1564);
    outputs(1674) <= not(layer0_outputs(1557));
    outputs(1675) <= (layer0_outputs(1268)) and not (layer0_outputs(1947));
    outputs(1676) <= not(layer0_outputs(480));
    outputs(1677) <= (layer0_outputs(129)) and (layer0_outputs(164));
    outputs(1678) <= not(layer0_outputs(2075));
    outputs(1679) <= layer0_outputs(14);
    outputs(1680) <= layer0_outputs(2003);
    outputs(1681) <= layer0_outputs(1327);
    outputs(1682) <= not(layer0_outputs(1266)) or (layer0_outputs(1122));
    outputs(1683) <= not((layer0_outputs(752)) or (layer0_outputs(1188)));
    outputs(1684) <= not(layer0_outputs(1412)) or (layer0_outputs(2356));
    outputs(1685) <= not((layer0_outputs(142)) xor (layer0_outputs(2405)));
    outputs(1686) <= not(layer0_outputs(1057));
    outputs(1687) <= not(layer0_outputs(1341));
    outputs(1688) <= (layer0_outputs(893)) and not (layer0_outputs(1985));
    outputs(1689) <= (layer0_outputs(1450)) and not (layer0_outputs(1243));
    outputs(1690) <= not(layer0_outputs(2513));
    outputs(1691) <= (layer0_outputs(123)) and not (layer0_outputs(924));
    outputs(1692) <= not((layer0_outputs(1972)) xor (layer0_outputs(1692)));
    outputs(1693) <= (layer0_outputs(2486)) and not (layer0_outputs(2072));
    outputs(1694) <= layer0_outputs(785);
    outputs(1695) <= not(layer0_outputs(924)) or (layer0_outputs(2165));
    outputs(1696) <= not((layer0_outputs(1028)) and (layer0_outputs(2317)));
    outputs(1697) <= not(layer0_outputs(557));
    outputs(1698) <= (layer0_outputs(1743)) and (layer0_outputs(1804));
    outputs(1699) <= layer0_outputs(973);
    outputs(1700) <= not(layer0_outputs(1025)) or (layer0_outputs(704));
    outputs(1701) <= layer0_outputs(722);
    outputs(1702) <= (layer0_outputs(286)) xor (layer0_outputs(1588));
    outputs(1703) <= layer0_outputs(1446);
    outputs(1704) <= not(layer0_outputs(260));
    outputs(1705) <= not((layer0_outputs(2346)) xor (layer0_outputs(1399)));
    outputs(1706) <= not(layer0_outputs(558));
    outputs(1707) <= (layer0_outputs(1178)) or (layer0_outputs(1067));
    outputs(1708) <= not(layer0_outputs(387));
    outputs(1709) <= not(layer0_outputs(2133));
    outputs(1710) <= (layer0_outputs(646)) and not (layer0_outputs(1948));
    outputs(1711) <= not(layer0_outputs(720));
    outputs(1712) <= (layer0_outputs(2100)) and not (layer0_outputs(582));
    outputs(1713) <= (layer0_outputs(112)) and not (layer0_outputs(2315));
    outputs(1714) <= layer0_outputs(2209);
    outputs(1715) <= not((layer0_outputs(1234)) or (layer0_outputs(2465)));
    outputs(1716) <= layer0_outputs(1715);
    outputs(1717) <= (layer0_outputs(2320)) xor (layer0_outputs(352));
    outputs(1718) <= layer0_outputs(1404);
    outputs(1719) <= not(layer0_outputs(484));
    outputs(1720) <= not((layer0_outputs(1828)) and (layer0_outputs(636)));
    outputs(1721) <= not(layer0_outputs(575)) or (layer0_outputs(958));
    outputs(1722) <= layer0_outputs(1593);
    outputs(1723) <= not(layer0_outputs(225)) or (layer0_outputs(2266));
    outputs(1724) <= not((layer0_outputs(790)) or (layer0_outputs(659)));
    outputs(1725) <= (layer0_outputs(13)) and not (layer0_outputs(638));
    outputs(1726) <= layer0_outputs(1706);
    outputs(1727) <= not((layer0_outputs(458)) xor (layer0_outputs(978)));
    outputs(1728) <= not((layer0_outputs(1643)) or (layer0_outputs(2067)));
    outputs(1729) <= not((layer0_outputs(772)) or (layer0_outputs(2168)));
    outputs(1730) <= not((layer0_outputs(288)) and (layer0_outputs(1910)));
    outputs(1731) <= not(layer0_outputs(928));
    outputs(1732) <= (layer0_outputs(506)) and (layer0_outputs(2332));
    outputs(1733) <= not(layer0_outputs(2352));
    outputs(1734) <= (layer0_outputs(808)) or (layer0_outputs(400));
    outputs(1735) <= (layer0_outputs(2559)) xor (layer0_outputs(1697));
    outputs(1736) <= (layer0_outputs(1398)) xor (layer0_outputs(1294));
    outputs(1737) <= layer0_outputs(1696);
    outputs(1738) <= (layer0_outputs(703)) xor (layer0_outputs(420));
    outputs(1739) <= not((layer0_outputs(1058)) and (layer0_outputs(2464)));
    outputs(1740) <= (layer0_outputs(1331)) and not (layer0_outputs(1162));
    outputs(1741) <= not(layer0_outputs(90));
    outputs(1742) <= not((layer0_outputs(1590)) or (layer0_outputs(1809)));
    outputs(1743) <= not(layer0_outputs(163));
    outputs(1744) <= not((layer0_outputs(2153)) or (layer0_outputs(2184)));
    outputs(1745) <= not(layer0_outputs(860));
    outputs(1746) <= (layer0_outputs(202)) and not (layer0_outputs(533));
    outputs(1747) <= not(layer0_outputs(441)) or (layer0_outputs(2406));
    outputs(1748) <= (layer0_outputs(34)) xor (layer0_outputs(832));
    outputs(1749) <= (layer0_outputs(1900)) and (layer0_outputs(1510));
    outputs(1750) <= (layer0_outputs(1805)) and not (layer0_outputs(1098));
    outputs(1751) <= layer0_outputs(1433);
    outputs(1752) <= not(layer0_outputs(1977));
    outputs(1753) <= not(layer0_outputs(445)) or (layer0_outputs(712));
    outputs(1754) <= not((layer0_outputs(258)) or (layer0_outputs(2120)));
    outputs(1755) <= layer0_outputs(2544);
    outputs(1756) <= (layer0_outputs(315)) and (layer0_outputs(995));
    outputs(1757) <= not(layer0_outputs(99)) or (layer0_outputs(1126));
    outputs(1758) <= (layer0_outputs(1059)) and not (layer0_outputs(1820));
    outputs(1759) <= layer0_outputs(2269);
    outputs(1760) <= not(layer0_outputs(2085)) or (layer0_outputs(310));
    outputs(1761) <= not((layer0_outputs(2430)) and (layer0_outputs(252)));
    outputs(1762) <= not(layer0_outputs(1834)) or (layer0_outputs(1061));
    outputs(1763) <= not(layer0_outputs(1040));
    outputs(1764) <= layer0_outputs(705);
    outputs(1765) <= not((layer0_outputs(891)) or (layer0_outputs(2227)));
    outputs(1766) <= (layer0_outputs(1896)) and not (layer0_outputs(1748));
    outputs(1767) <= not(layer0_outputs(1660));
    outputs(1768) <= not((layer0_outputs(1781)) xor (layer0_outputs(21)));
    outputs(1769) <= not(layer0_outputs(2146));
    outputs(1770) <= (layer0_outputs(1356)) and (layer0_outputs(640));
    outputs(1771) <= (layer0_outputs(1029)) xor (layer0_outputs(1581));
    outputs(1772) <= not(layer0_outputs(2507));
    outputs(1773) <= (layer0_outputs(169)) xor (layer0_outputs(1790));
    outputs(1774) <= layer0_outputs(1530);
    outputs(1775) <= layer0_outputs(2152);
    outputs(1776) <= (layer0_outputs(925)) and not (layer0_outputs(2418));
    outputs(1777) <= (layer0_outputs(390)) and (layer0_outputs(1687));
    outputs(1778) <= (layer0_outputs(2415)) xor (layer0_outputs(2318));
    outputs(1779) <= not(layer0_outputs(2423));
    outputs(1780) <= (layer0_outputs(1263)) and (layer0_outputs(1136));
    outputs(1781) <= (layer0_outputs(757)) and not (layer0_outputs(2249));
    outputs(1782) <= not((layer0_outputs(1207)) or (layer0_outputs(766)));
    outputs(1783) <= not((layer0_outputs(150)) or (layer0_outputs(342)));
    outputs(1784) <= (layer0_outputs(433)) and not (layer0_outputs(1202));
    outputs(1785) <= (layer0_outputs(2327)) and not (layer0_outputs(1174));
    outputs(1786) <= (layer0_outputs(1476)) and not (layer0_outputs(1044));
    outputs(1787) <= (layer0_outputs(801)) and (layer0_outputs(1541));
    outputs(1788) <= (layer0_outputs(2078)) and not (layer0_outputs(1948));
    outputs(1789) <= layer0_outputs(2100);
    outputs(1790) <= not((layer0_outputs(1905)) and (layer0_outputs(95)));
    outputs(1791) <= (layer0_outputs(1881)) and not (layer0_outputs(1855));
    outputs(1792) <= not((layer0_outputs(2307)) and (layer0_outputs(98)));
    outputs(1793) <= not(layer0_outputs(255));
    outputs(1794) <= (layer0_outputs(1666)) xor (layer0_outputs(1932));
    outputs(1795) <= not((layer0_outputs(2413)) xor (layer0_outputs(314)));
    outputs(1796) <= (layer0_outputs(1165)) and not (layer0_outputs(1530));
    outputs(1797) <= (layer0_outputs(1272)) and not (layer0_outputs(1331));
    outputs(1798) <= not(layer0_outputs(1989)) or (layer0_outputs(912));
    outputs(1799) <= layer0_outputs(2384);
    outputs(1800) <= (layer0_outputs(715)) and not (layer0_outputs(1064));
    outputs(1801) <= (layer0_outputs(118)) xor (layer0_outputs(1079));
    outputs(1802) <= (layer0_outputs(138)) and (layer0_outputs(1991));
    outputs(1803) <= not(layer0_outputs(276));
    outputs(1804) <= (layer0_outputs(742)) xor (layer0_outputs(934));
    outputs(1805) <= layer0_outputs(1596);
    outputs(1806) <= not(layer0_outputs(1895));
    outputs(1807) <= not((layer0_outputs(488)) or (layer0_outputs(1397)));
    outputs(1808) <= not((layer0_outputs(1208)) xor (layer0_outputs(46)));
    outputs(1809) <= layer0_outputs(2260);
    outputs(1810) <= not((layer0_outputs(1016)) or (layer0_outputs(1507)));
    outputs(1811) <= '1';
    outputs(1812) <= not(layer0_outputs(2002)) or (layer0_outputs(153));
    outputs(1813) <= not((layer0_outputs(1722)) or (layer0_outputs(686)));
    outputs(1814) <= not((layer0_outputs(1044)) or (layer0_outputs(783)));
    outputs(1815) <= layer0_outputs(2270);
    outputs(1816) <= not(layer0_outputs(2343)) or (layer0_outputs(1452));
    outputs(1817) <= not(layer0_outputs(656));
    outputs(1818) <= layer0_outputs(900);
    outputs(1819) <= (layer0_outputs(2129)) xor (layer0_outputs(1061));
    outputs(1820) <= not(layer0_outputs(386));
    outputs(1821) <= (layer0_outputs(1103)) and not (layer0_outputs(1569));
    outputs(1822) <= (layer0_outputs(170)) and (layer0_outputs(896));
    outputs(1823) <= (layer0_outputs(893)) xor (layer0_outputs(1518));
    outputs(1824) <= not(layer0_outputs(248));
    outputs(1825) <= not((layer0_outputs(630)) or (layer0_outputs(2277)));
    outputs(1826) <= (layer0_outputs(1759)) and not (layer0_outputs(1899));
    outputs(1827) <= not((layer0_outputs(1591)) or (layer0_outputs(989)));
    outputs(1828) <= not(layer0_outputs(490));
    outputs(1829) <= (layer0_outputs(1726)) and not (layer0_outputs(1116));
    outputs(1830) <= not((layer0_outputs(1529)) xor (layer0_outputs(841)));
    outputs(1831) <= not(layer0_outputs(639));
    outputs(1832) <= (layer0_outputs(1732)) and not (layer0_outputs(2410));
    outputs(1833) <= not(layer0_outputs(2316));
    outputs(1834) <= (layer0_outputs(1438)) and not (layer0_outputs(1217));
    outputs(1835) <= (layer0_outputs(1416)) xor (layer0_outputs(1554));
    outputs(1836) <= layer0_outputs(247);
    outputs(1837) <= not(layer0_outputs(314));
    outputs(1838) <= not((layer0_outputs(1142)) xor (layer0_outputs(2098)));
    outputs(1839) <= (layer0_outputs(837)) xor (layer0_outputs(139));
    outputs(1840) <= (layer0_outputs(976)) and (layer0_outputs(1042));
    outputs(1841) <= not(layer0_outputs(901));
    outputs(1842) <= not(layer0_outputs(2470));
    outputs(1843) <= not((layer0_outputs(685)) and (layer0_outputs(1779)));
    outputs(1844) <= not(layer0_outputs(1297));
    outputs(1845) <= (layer0_outputs(1286)) xor (layer0_outputs(774));
    outputs(1846) <= not(layer0_outputs(960)) or (layer0_outputs(1688));
    outputs(1847) <= '0';
    outputs(1848) <= not(layer0_outputs(357));
    outputs(1849) <= not(layer0_outputs(1031));
    outputs(1850) <= not((layer0_outputs(1035)) or (layer0_outputs(1037)));
    outputs(1851) <= not((layer0_outputs(749)) xor (layer0_outputs(1389)));
    outputs(1852) <= (layer0_outputs(2096)) xor (layer0_outputs(1681));
    outputs(1853) <= not((layer0_outputs(1785)) or (layer0_outputs(1002)));
    outputs(1854) <= not((layer0_outputs(2343)) xor (layer0_outputs(1602)));
    outputs(1855) <= (layer0_outputs(2090)) xor (layer0_outputs(1151));
    outputs(1856) <= (layer0_outputs(851)) and not (layer0_outputs(166));
    outputs(1857) <= (layer0_outputs(187)) xor (layer0_outputs(1421));
    outputs(1858) <= not(layer0_outputs(2052)) or (layer0_outputs(230));
    outputs(1859) <= not(layer0_outputs(73));
    outputs(1860) <= layer0_outputs(2483);
    outputs(1861) <= layer0_outputs(2463);
    outputs(1862) <= (layer0_outputs(1794)) and not (layer0_outputs(1831));
    outputs(1863) <= not(layer0_outputs(2142));
    outputs(1864) <= not((layer0_outputs(1121)) or (layer0_outputs(83)));
    outputs(1865) <= (layer0_outputs(1946)) and not (layer0_outputs(767));
    outputs(1866) <= layer0_outputs(1119);
    outputs(1867) <= not((layer0_outputs(229)) or (layer0_outputs(1060)));
    outputs(1868) <= not(layer0_outputs(1984));
    outputs(1869) <= (layer0_outputs(2263)) and not (layer0_outputs(935));
    outputs(1870) <= not(layer0_outputs(298));
    outputs(1871) <= not((layer0_outputs(207)) or (layer0_outputs(810)));
    outputs(1872) <= not(layer0_outputs(642));
    outputs(1873) <= not(layer0_outputs(126));
    outputs(1874) <= (layer0_outputs(1408)) and (layer0_outputs(4));
    outputs(1875) <= (layer0_outputs(1636)) and not (layer0_outputs(410));
    outputs(1876) <= not((layer0_outputs(1936)) xor (layer0_outputs(2288)));
    outputs(1877) <= layer0_outputs(573);
    outputs(1878) <= (layer0_outputs(316)) xor (layer0_outputs(0));
    outputs(1879) <= (layer0_outputs(621)) and not (layer0_outputs(933));
    outputs(1880) <= (layer0_outputs(557)) and not (layer0_outputs(1622));
    outputs(1881) <= not(layer0_outputs(2550)) or (layer0_outputs(1853));
    outputs(1882) <= (layer0_outputs(2448)) and (layer0_outputs(1081));
    outputs(1883) <= not(layer0_outputs(53));
    outputs(1884) <= layer0_outputs(1200);
    outputs(1885) <= not((layer0_outputs(800)) or (layer0_outputs(881)));
    outputs(1886) <= layer0_outputs(872);
    outputs(1887) <= not(layer0_outputs(1456));
    outputs(1888) <= (layer0_outputs(2131)) xor (layer0_outputs(2475));
    outputs(1889) <= (layer0_outputs(1209)) xor (layer0_outputs(2098));
    outputs(1890) <= (layer0_outputs(1499)) and not (layer0_outputs(1539));
    outputs(1891) <= not((layer0_outputs(878)) xor (layer0_outputs(523)));
    outputs(1892) <= (layer0_outputs(2193)) xor (layer0_outputs(970));
    outputs(1893) <= layer0_outputs(803);
    outputs(1894) <= layer0_outputs(1034);
    outputs(1895) <= not((layer0_outputs(1733)) and (layer0_outputs(937)));
    outputs(1896) <= not(layer0_outputs(981));
    outputs(1897) <= (layer0_outputs(2184)) xor (layer0_outputs(2443));
    outputs(1898) <= (layer0_outputs(495)) xor (layer0_outputs(1642));
    outputs(1899) <= (layer0_outputs(191)) and not (layer0_outputs(1496));
    outputs(1900) <= not(layer0_outputs(87));
    outputs(1901) <= not(layer0_outputs(26));
    outputs(1902) <= (layer0_outputs(1841)) and not (layer0_outputs(830));
    outputs(1903) <= not(layer0_outputs(696)) or (layer0_outputs(2340));
    outputs(1904) <= layer0_outputs(745);
    outputs(1905) <= (layer0_outputs(2181)) and (layer0_outputs(747));
    outputs(1906) <= not((layer0_outputs(2367)) and (layer0_outputs(1078)));
    outputs(1907) <= layer0_outputs(1525);
    outputs(1908) <= not(layer0_outputs(882));
    outputs(1909) <= not(layer0_outputs(174));
    outputs(1910) <= layer0_outputs(349);
    outputs(1911) <= (layer0_outputs(2238)) or (layer0_outputs(1099));
    outputs(1912) <= layer0_outputs(914);
    outputs(1913) <= layer0_outputs(1561);
    outputs(1914) <= not(layer0_outputs(897));
    outputs(1915) <= layer0_outputs(2534);
    outputs(1916) <= not(layer0_outputs(1581));
    outputs(1917) <= not((layer0_outputs(956)) xor (layer0_outputs(256)));
    outputs(1918) <= not(layer0_outputs(1507));
    outputs(1919) <= not(layer0_outputs(897));
    outputs(1920) <= layer0_outputs(1771);
    outputs(1921) <= not((layer0_outputs(2335)) or (layer0_outputs(692)));
    outputs(1922) <= not((layer0_outputs(350)) or (layer0_outputs(1090)));
    outputs(1923) <= not((layer0_outputs(1503)) or (layer0_outputs(2348)));
    outputs(1924) <= not((layer0_outputs(114)) xor (layer0_outputs(156)));
    outputs(1925) <= (layer0_outputs(847)) or (layer0_outputs(1858));
    outputs(1926) <= layer0_outputs(2039);
    outputs(1927) <= layer0_outputs(1666);
    outputs(1928) <= not((layer0_outputs(2480)) and (layer0_outputs(1078)));
    outputs(1929) <= (layer0_outputs(318)) or (layer0_outputs(681));
    outputs(1930) <= not((layer0_outputs(1252)) or (layer0_outputs(831)));
    outputs(1931) <= (layer0_outputs(2148)) and not (layer0_outputs(1222));
    outputs(1932) <= not(layer0_outputs(2431));
    outputs(1933) <= not(layer0_outputs(693));
    outputs(1934) <= not(layer0_outputs(1856));
    outputs(1935) <= (layer0_outputs(1523)) xor (layer0_outputs(931));
    outputs(1936) <= (layer0_outputs(611)) or (layer0_outputs(327));
    outputs(1937) <= layer0_outputs(688);
    outputs(1938) <= not(layer0_outputs(2477));
    outputs(1939) <= layer0_outputs(303);
    outputs(1940) <= not((layer0_outputs(1112)) or (layer0_outputs(1309)));
    outputs(1941) <= layer0_outputs(204);
    outputs(1942) <= not((layer0_outputs(400)) xor (layer0_outputs(797)));
    outputs(1943) <= not(layer0_outputs(594));
    outputs(1944) <= not(layer0_outputs(748));
    outputs(1945) <= not(layer0_outputs(1931));
    outputs(1946) <= not(layer0_outputs(1138));
    outputs(1947) <= layer0_outputs(2178);
    outputs(1948) <= (layer0_outputs(137)) and not (layer0_outputs(52));
    outputs(1949) <= not(layer0_outputs(2239));
    outputs(1950) <= not((layer0_outputs(1678)) xor (layer0_outputs(1799)));
    outputs(1951) <= not(layer0_outputs(1959));
    outputs(1952) <= not(layer0_outputs(102));
    outputs(1953) <= not(layer0_outputs(1411));
    outputs(1954) <= not(layer0_outputs(2390));
    outputs(1955) <= not(layer0_outputs(887)) or (layer0_outputs(2507));
    outputs(1956) <= not((layer0_outputs(55)) or (layer0_outputs(18)));
    outputs(1957) <= (layer0_outputs(618)) and (layer0_outputs(1974));
    outputs(1958) <= not(layer0_outputs(1980));
    outputs(1959) <= not(layer0_outputs(1150));
    outputs(1960) <= not(layer0_outputs(2198));
    outputs(1961) <= (layer0_outputs(1946)) and (layer0_outputs(2176));
    outputs(1962) <= not((layer0_outputs(155)) xor (layer0_outputs(845)));
    outputs(1963) <= not(layer0_outputs(1654));
    outputs(1964) <= (layer0_outputs(1320)) xor (layer0_outputs(953));
    outputs(1965) <= (layer0_outputs(1108)) and not (layer0_outputs(2225));
    outputs(1966) <= (layer0_outputs(2295)) and not (layer0_outputs(2276));
    outputs(1967) <= not((layer0_outputs(1198)) xor (layer0_outputs(738)));
    outputs(1968) <= (layer0_outputs(1190)) and (layer0_outputs(1634));
    outputs(1969) <= not(layer0_outputs(555));
    outputs(1970) <= not(layer0_outputs(2014));
    outputs(1971) <= layer0_outputs(524);
    outputs(1972) <= (layer0_outputs(1091)) xor (layer0_outputs(692));
    outputs(1973) <= layer0_outputs(698);
    outputs(1974) <= (layer0_outputs(1436)) and not (layer0_outputs(475));
    outputs(1975) <= layer0_outputs(698);
    outputs(1976) <= layer0_outputs(430);
    outputs(1977) <= layer0_outputs(1394);
    outputs(1978) <= layer0_outputs(1903);
    outputs(1979) <= not(layer0_outputs(2113));
    outputs(1980) <= (layer0_outputs(1766)) xor (layer0_outputs(626));
    outputs(1981) <= (layer0_outputs(2055)) and not (layer0_outputs(24));
    outputs(1982) <= (layer0_outputs(1702)) xor (layer0_outputs(1852));
    outputs(1983) <= (layer0_outputs(2445)) and not (layer0_outputs(789));
    outputs(1984) <= not(layer0_outputs(739));
    outputs(1985) <= not(layer0_outputs(2452));
    outputs(1986) <= (layer0_outputs(1625)) and not (layer0_outputs(1233));
    outputs(1987) <= (layer0_outputs(282)) or (layer0_outputs(714));
    outputs(1988) <= layer0_outputs(1467);
    outputs(1989) <= not(layer0_outputs(332));
    outputs(1990) <= (layer0_outputs(1408)) and not (layer0_outputs(2312));
    outputs(1991) <= not((layer0_outputs(2341)) xor (layer0_outputs(218)));
    outputs(1992) <= not(layer0_outputs(1651));
    outputs(1993) <= (layer0_outputs(1907)) and not (layer0_outputs(1950));
    outputs(1994) <= not(layer0_outputs(1859)) or (layer0_outputs(585));
    outputs(1995) <= (layer0_outputs(1071)) and not (layer0_outputs(1669));
    outputs(1996) <= (layer0_outputs(982)) xor (layer0_outputs(588));
    outputs(1997) <= layer0_outputs(42);
    outputs(1998) <= not(layer0_outputs(2284));
    outputs(1999) <= not(layer0_outputs(2239)) or (layer0_outputs(115));
    outputs(2000) <= not((layer0_outputs(1113)) or (layer0_outputs(2398)));
    outputs(2001) <= not((layer0_outputs(2095)) xor (layer0_outputs(584)));
    outputs(2002) <= not((layer0_outputs(1545)) or (layer0_outputs(110)));
    outputs(2003) <= not(layer0_outputs(818));
    outputs(2004) <= not((layer0_outputs(1009)) xor (layer0_outputs(2404)));
    outputs(2005) <= (layer0_outputs(1865)) and not (layer0_outputs(402));
    outputs(2006) <= (layer0_outputs(1474)) and not (layer0_outputs(1549));
    outputs(2007) <= (layer0_outputs(2144)) and (layer0_outputs(578));
    outputs(2008) <= (layer0_outputs(794)) and not (layer0_outputs(486));
    outputs(2009) <= layer0_outputs(2432);
    outputs(2010) <= layer0_outputs(2490);
    outputs(2011) <= not((layer0_outputs(1888)) or (layer0_outputs(1693)));
    outputs(2012) <= not((layer0_outputs(2034)) or (layer0_outputs(1565)));
    outputs(2013) <= (layer0_outputs(1193)) and (layer0_outputs(38));
    outputs(2014) <= not((layer0_outputs(670)) and (layer0_outputs(905)));
    outputs(2015) <= not((layer0_outputs(1807)) or (layer0_outputs(459)));
    outputs(2016) <= (layer0_outputs(808)) xor (layer0_outputs(1204));
    outputs(2017) <= (layer0_outputs(967)) and (layer0_outputs(1649));
    outputs(2018) <= layer0_outputs(2365);
    outputs(2019) <= layer0_outputs(1567);
    outputs(2020) <= layer0_outputs(167);
    outputs(2021) <= not(layer0_outputs(249));
    outputs(2022) <= not(layer0_outputs(320));
    outputs(2023) <= (layer0_outputs(1027)) or (layer0_outputs(2355));
    outputs(2024) <= not(layer0_outputs(1123)) or (layer0_outputs(1148));
    outputs(2025) <= layer0_outputs(1854);
    outputs(2026) <= not(layer0_outputs(380)) or (layer0_outputs(1897));
    outputs(2027) <= layer0_outputs(44);
    outputs(2028) <= not(layer0_outputs(776));
    outputs(2029) <= not(layer0_outputs(2230));
    outputs(2030) <= (layer0_outputs(1328)) xor (layer0_outputs(1090));
    outputs(2031) <= not((layer0_outputs(1659)) xor (layer0_outputs(1453)));
    outputs(2032) <= not((layer0_outputs(1171)) or (layer0_outputs(321)));
    outputs(2033) <= not((layer0_outputs(1916)) or (layer0_outputs(125)));
    outputs(2034) <= not(layer0_outputs(397)) or (layer0_outputs(1228));
    outputs(2035) <= (layer0_outputs(1291)) and (layer0_outputs(2087));
    outputs(2036) <= (layer0_outputs(372)) xor (layer0_outputs(1145));
    outputs(2037) <= layer0_outputs(2454);
    outputs(2038) <= not(layer0_outputs(2073));
    outputs(2039) <= not((layer0_outputs(769)) or (layer0_outputs(2335)));
    outputs(2040) <= layer0_outputs(29);
    outputs(2041) <= not(layer0_outputs(741));
    outputs(2042) <= layer0_outputs(2022);
    outputs(2043) <= not(layer0_outputs(2065));
    outputs(2044) <= (layer0_outputs(823)) and (layer0_outputs(423));
    outputs(2045) <= (layer0_outputs(1760)) or (layer0_outputs(1988));
    outputs(2046) <= not(layer0_outputs(2088));
    outputs(2047) <= (layer0_outputs(1156)) and not (layer0_outputs(1661));
    outputs(2048) <= not((layer0_outputs(1406)) or (layer0_outputs(1425)));
    outputs(2049) <= layer0_outputs(2472);
    outputs(2050) <= not((layer0_outputs(2063)) and (layer0_outputs(2508)));
    outputs(2051) <= (layer0_outputs(719)) or (layer0_outputs(2500));
    outputs(2052) <= not(layer0_outputs(2538));
    outputs(2053) <= layer0_outputs(925);
    outputs(2054) <= not(layer0_outputs(1555));
    outputs(2055) <= not((layer0_outputs(1313)) and (layer0_outputs(2511)));
    outputs(2056) <= (layer0_outputs(1624)) and (layer0_outputs(2529));
    outputs(2057) <= (layer0_outputs(2275)) and (layer0_outputs(1428));
    outputs(2058) <= not(layer0_outputs(2374));
    outputs(2059) <= not(layer0_outputs(578));
    outputs(2060) <= not(layer0_outputs(1169));
    outputs(2061) <= layer0_outputs(1884);
    outputs(2062) <= not((layer0_outputs(1925)) xor (layer0_outputs(1380)));
    outputs(2063) <= (layer0_outputs(1974)) and (layer0_outputs(2257));
    outputs(2064) <= layer0_outputs(1010);
    outputs(2065) <= not(layer0_outputs(910));
    outputs(2066) <= (layer0_outputs(689)) xor (layer0_outputs(477));
    outputs(2067) <= (layer0_outputs(1716)) and not (layer0_outputs(630));
    outputs(2068) <= not(layer0_outputs(1041)) or (layer0_outputs(2482));
    outputs(2069) <= not(layer0_outputs(47)) or (layer0_outputs(1163));
    outputs(2070) <= not((layer0_outputs(857)) or (layer0_outputs(288)));
    outputs(2071) <= not((layer0_outputs(915)) xor (layer0_outputs(2328)));
    outputs(2072) <= not(layer0_outputs(485)) or (layer0_outputs(1244));
    outputs(2073) <= (layer0_outputs(812)) and not (layer0_outputs(1275));
    outputs(2074) <= not(layer0_outputs(148));
    outputs(2075) <= (layer0_outputs(176)) and not (layer0_outputs(711));
    outputs(2076) <= (layer0_outputs(743)) and not (layer0_outputs(1739));
    outputs(2077) <= (layer0_outputs(610)) and not (layer0_outputs(1190));
    outputs(2078) <= layer0_outputs(1966);
    outputs(2079) <= not(layer0_outputs(1026));
    outputs(2080) <= layer0_outputs(614);
    outputs(2081) <= not((layer0_outputs(2515)) xor (layer0_outputs(2471)));
    outputs(2082) <= not(layer0_outputs(1797));
    outputs(2083) <= (layer0_outputs(515)) xor (layer0_outputs(1322));
    outputs(2084) <= layer0_outputs(522);
    outputs(2085) <= (layer0_outputs(1223)) and not (layer0_outputs(131));
    outputs(2086) <= not(layer0_outputs(1537));
    outputs(2087) <= not((layer0_outputs(182)) or (layer0_outputs(196)));
    outputs(2088) <= not(layer0_outputs(39));
    outputs(2089) <= not(layer0_outputs(2535));
    outputs(2090) <= not((layer0_outputs(2351)) xor (layer0_outputs(2359)));
    outputs(2091) <= not((layer0_outputs(862)) or (layer0_outputs(688)));
    outputs(2092) <= not((layer0_outputs(2383)) and (layer0_outputs(992)));
    outputs(2093) <= not((layer0_outputs(582)) or (layer0_outputs(623)));
    outputs(2094) <= (layer0_outputs(2265)) and not (layer0_outputs(1640));
    outputs(2095) <= layer0_outputs(740);
    outputs(2096) <= layer0_outputs(2378);
    outputs(2097) <= (layer0_outputs(2342)) and (layer0_outputs(1545));
    outputs(2098) <= (layer0_outputs(2412)) xor (layer0_outputs(2160));
    outputs(2099) <= not(layer0_outputs(1177));
    outputs(2100) <= not((layer0_outputs(2091)) xor (layer0_outputs(850)));
    outputs(2101) <= layer0_outputs(1928);
    outputs(2102) <= not((layer0_outputs(2046)) or (layer0_outputs(1487)));
    outputs(2103) <= (layer0_outputs(171)) xor (layer0_outputs(1757));
    outputs(2104) <= not(layer0_outputs(371));
    outputs(2105) <= not(layer0_outputs(2374));
    outputs(2106) <= (layer0_outputs(1707)) and (layer0_outputs(778));
    outputs(2107) <= not((layer0_outputs(487)) xor (layer0_outputs(163)));
    outputs(2108) <= not((layer0_outputs(377)) xor (layer0_outputs(291)));
    outputs(2109) <= (layer0_outputs(952)) and not (layer0_outputs(1470));
    outputs(2110) <= (layer0_outputs(683)) and not (layer0_outputs(2454));
    outputs(2111) <= not(layer0_outputs(181)) or (layer0_outputs(2345));
    outputs(2112) <= layer0_outputs(8);
    outputs(2113) <= not(layer0_outputs(712));
    outputs(2114) <= layer0_outputs(1650);
    outputs(2115) <= not((layer0_outputs(126)) xor (layer0_outputs(496)));
    outputs(2116) <= layer0_outputs(307);
    outputs(2117) <= not((layer0_outputs(753)) xor (layer0_outputs(1431)));
    outputs(2118) <= not(layer0_outputs(2112));
    outputs(2119) <= not((layer0_outputs(374)) xor (layer0_outputs(1407)));
    outputs(2120) <= not(layer0_outputs(982)) or (layer0_outputs(1321));
    outputs(2121) <= not((layer0_outputs(583)) xor (layer0_outputs(2037)));
    outputs(2122) <= (layer0_outputs(397)) and (layer0_outputs(360));
    outputs(2123) <= not(layer0_outputs(2512));
    outputs(2124) <= (layer0_outputs(1251)) and not (layer0_outputs(2118));
    outputs(2125) <= (layer0_outputs(2553)) and (layer0_outputs(1843));
    outputs(2126) <= not(layer0_outputs(1825)) or (layer0_outputs(789));
    outputs(2127) <= (layer0_outputs(2154)) and (layer0_outputs(1328));
    outputs(2128) <= not(layer0_outputs(1668));
    outputs(2129) <= not((layer0_outputs(1069)) xor (layer0_outputs(1492)));
    outputs(2130) <= not((layer0_outputs(1460)) xor (layer0_outputs(1618)));
    outputs(2131) <= (layer0_outputs(1978)) and not (layer0_outputs(490));
    outputs(2132) <= not((layer0_outputs(1730)) or (layer0_outputs(451)));
    outputs(2133) <= not((layer0_outputs(2229)) xor (layer0_outputs(2483)));
    outputs(2134) <= (layer0_outputs(1659)) and not (layer0_outputs(271));
    outputs(2135) <= layer0_outputs(1273);
    outputs(2136) <= layer0_outputs(1704);
    outputs(2137) <= not(layer0_outputs(744)) or (layer0_outputs(23));
    outputs(2138) <= (layer0_outputs(143)) xor (layer0_outputs(600));
    outputs(2139) <= not(layer0_outputs(1569));
    outputs(2140) <= layer0_outputs(733);
    outputs(2141) <= (layer0_outputs(2457)) and not (layer0_outputs(1528));
    outputs(2142) <= (layer0_outputs(1920)) and (layer0_outputs(552));
    outputs(2143) <= not(layer0_outputs(966));
    outputs(2144) <= (layer0_outputs(1749)) and (layer0_outputs(308));
    outputs(2145) <= not((layer0_outputs(1868)) or (layer0_outputs(2011)));
    outputs(2146) <= not(layer0_outputs(364));
    outputs(2147) <= not(layer0_outputs(164));
    outputs(2148) <= not(layer0_outputs(2381));
    outputs(2149) <= not(layer0_outputs(1720));
    outputs(2150) <= layer0_outputs(894);
    outputs(2151) <= not(layer0_outputs(422));
    outputs(2152) <= (layer0_outputs(943)) and not (layer0_outputs(2037));
    outputs(2153) <= not(layer0_outputs(1309));
    outputs(2154) <= not((layer0_outputs(1259)) xor (layer0_outputs(1717)));
    outputs(2155) <= (layer0_outputs(2023)) and not (layer0_outputs(2282));
    outputs(2156) <= not(layer0_outputs(999));
    outputs(2157) <= not((layer0_outputs(751)) or (layer0_outputs(1308)));
    outputs(2158) <= layer0_outputs(798);
    outputs(2159) <= not((layer0_outputs(689)) xor (layer0_outputs(1458)));
    outputs(2160) <= (layer0_outputs(829)) and not (layer0_outputs(1644));
    outputs(2161) <= layer0_outputs(1811);
    outputs(2162) <= not((layer0_outputs(1014)) and (layer0_outputs(1041)));
    outputs(2163) <= layer0_outputs(1131);
    outputs(2164) <= not(layer0_outputs(1806));
    outputs(2165) <= (layer0_outputs(786)) and not (layer0_outputs(428));
    outputs(2166) <= layer0_outputs(2268);
    outputs(2167) <= not((layer0_outputs(1911)) or (layer0_outputs(2418)));
    outputs(2168) <= not((layer0_outputs(823)) or (layer0_outputs(2050)));
    outputs(2169) <= (layer0_outputs(1694)) and not (layer0_outputs(658));
    outputs(2170) <= not((layer0_outputs(1937)) xor (layer0_outputs(2052)));
    outputs(2171) <= not(layer0_outputs(1969));
    outputs(2172) <= not((layer0_outputs(1531)) xor (layer0_outputs(1767)));
    outputs(2173) <= not(layer0_outputs(1371));
    outputs(2174) <= not(layer0_outputs(2369));
    outputs(2175) <= layer0_outputs(1887);
    outputs(2176) <= not((layer0_outputs(2478)) xor (layer0_outputs(824)));
    outputs(2177) <= not(layer0_outputs(2231));
    outputs(2178) <= not(layer0_outputs(1210));
    outputs(2179) <= (layer0_outputs(2106)) and (layer0_outputs(631));
    outputs(2180) <= layer0_outputs(2277);
    outputs(2181) <= not(layer0_outputs(476));
    outputs(2182) <= (layer0_outputs(2476)) and (layer0_outputs(1367));
    outputs(2183) <= layer0_outputs(468);
    outputs(2184) <= layer0_outputs(152);
    outputs(2185) <= (layer0_outputs(267)) and (layer0_outputs(1816));
    outputs(2186) <= (layer0_outputs(1223)) xor (layer0_outputs(1322));
    outputs(2187) <= not(layer0_outputs(1280));
    outputs(2188) <= (layer0_outputs(817)) and not (layer0_outputs(1118));
    outputs(2189) <= not(layer0_outputs(1980));
    outputs(2190) <= (layer0_outputs(2104)) and not (layer0_outputs(919));
    outputs(2191) <= not(layer0_outputs(837));
    outputs(2192) <= not((layer0_outputs(1595)) xor (layer0_outputs(1203)));
    outputs(2193) <= (layer0_outputs(82)) xor (layer0_outputs(1437));
    outputs(2194) <= (layer0_outputs(68)) xor (layer0_outputs(2030));
    outputs(2195) <= not(layer0_outputs(832)) or (layer0_outputs(460));
    outputs(2196) <= (layer0_outputs(987)) and not (layer0_outputs(237));
    outputs(2197) <= not(layer0_outputs(2300)) or (layer0_outputs(159));
    outputs(2198) <= (layer0_outputs(1582)) and not (layer0_outputs(1036));
    outputs(2199) <= not((layer0_outputs(1257)) xor (layer0_outputs(1055)));
    outputs(2200) <= (layer0_outputs(1159)) and not (layer0_outputs(287));
    outputs(2201) <= (layer0_outputs(886)) and not (layer0_outputs(365));
    outputs(2202) <= not((layer0_outputs(1111)) xor (layer0_outputs(1849)));
    outputs(2203) <= not(layer0_outputs(1307)) or (layer0_outputs(918));
    outputs(2204) <= (layer0_outputs(1157)) and (layer0_outputs(1346));
    outputs(2205) <= (layer0_outputs(1262)) or (layer0_outputs(784));
    outputs(2206) <= (layer0_outputs(2208)) xor (layer0_outputs(1467));
    outputs(2207) <= layer0_outputs(782);
    outputs(2208) <= not((layer0_outputs(76)) xor (layer0_outputs(2287)));
    outputs(2209) <= (layer0_outputs(284)) and not (layer0_outputs(2420));
    outputs(2210) <= not((layer0_outputs(1191)) and (layer0_outputs(969)));
    outputs(2211) <= not((layer0_outputs(1777)) and (layer0_outputs(1652)));
    outputs(2212) <= not(layer0_outputs(208));
    outputs(2213) <= (layer0_outputs(173)) and not (layer0_outputs(1879));
    outputs(2214) <= (layer0_outputs(1971)) and (layer0_outputs(1146));
    outputs(2215) <= not(layer0_outputs(1345));
    outputs(2216) <= (layer0_outputs(1613)) xor (layer0_outputs(972));
    outputs(2217) <= not(layer0_outputs(2429));
    outputs(2218) <= not((layer0_outputs(406)) xor (layer0_outputs(1909)));
    outputs(2219) <= (layer0_outputs(1114)) and not (layer0_outputs(2245));
    outputs(2220) <= layer0_outputs(303);
    outputs(2221) <= not(layer0_outputs(2536));
    outputs(2222) <= (layer0_outputs(1570)) xor (layer0_outputs(2137));
    outputs(2223) <= (layer0_outputs(1986)) and not (layer0_outputs(2059));
    outputs(2224) <= (layer0_outputs(1691)) and not (layer0_outputs(1169));
    outputs(2225) <= not(layer0_outputs(1751));
    outputs(2226) <= (layer0_outputs(2097)) and not (layer0_outputs(691));
    outputs(2227) <= (layer0_outputs(435)) xor (layer0_outputs(1269));
    outputs(2228) <= (layer0_outputs(1746)) xor (layer0_outputs(2486));
    outputs(2229) <= not(layer0_outputs(840));
    outputs(2230) <= not(layer0_outputs(1341));
    outputs(2231) <= (layer0_outputs(1610)) or (layer0_outputs(1107));
    outputs(2232) <= not((layer0_outputs(2460)) or (layer0_outputs(2545)));
    outputs(2233) <= (layer0_outputs(1653)) and (layer0_outputs(1005));
    outputs(2234) <= (layer0_outputs(562)) xor (layer0_outputs(1743));
    outputs(2235) <= (layer0_outputs(1367)) and not (layer0_outputs(2327));
    outputs(2236) <= not(layer0_outputs(860));
    outputs(2237) <= not(layer0_outputs(447)) or (layer0_outputs(1635));
    outputs(2238) <= layer0_outputs(2283);
    outputs(2239) <= not(layer0_outputs(736));
    outputs(2240) <= not(layer0_outputs(1393));
    outputs(2241) <= not(layer0_outputs(1992));
    outputs(2242) <= not(layer0_outputs(1989));
    outputs(2243) <= (layer0_outputs(313)) and not (layer0_outputs(1627));
    outputs(2244) <= not(layer0_outputs(2274)) or (layer0_outputs(2082));
    outputs(2245) <= (layer0_outputs(338)) and (layer0_outputs(1230));
    outputs(2246) <= (layer0_outputs(137)) and not (layer0_outputs(529));
    outputs(2247) <= layer0_outputs(1429);
    outputs(2248) <= layer0_outputs(332);
    outputs(2249) <= not(layer0_outputs(984)) or (layer0_outputs(2385));
    outputs(2250) <= (layer0_outputs(1257)) and (layer0_outputs(1143));
    outputs(2251) <= not(layer0_outputs(709));
    outputs(2252) <= not(layer0_outputs(158));
    outputs(2253) <= not(layer0_outputs(89));
    outputs(2254) <= not((layer0_outputs(2125)) xor (layer0_outputs(2364)));
    outputs(2255) <= (layer0_outputs(2456)) and (layer0_outputs(1131));
    outputs(2256) <= layer0_outputs(1674);
    outputs(2257) <= not(layer0_outputs(1813)) or (layer0_outputs(917));
    outputs(2258) <= not(layer0_outputs(1782));
    outputs(2259) <= (layer0_outputs(2428)) and (layer0_outputs(1509));
    outputs(2260) <= not(layer0_outputs(2420));
    outputs(2261) <= not(layer0_outputs(102));
    outputs(2262) <= not((layer0_outputs(2466)) or (layer0_outputs(545)));
    outputs(2263) <= layer0_outputs(1196);
    outputs(2264) <= not((layer0_outputs(690)) xor (layer0_outputs(1664)));
    outputs(2265) <= layer0_outputs(1364);
    outputs(2266) <= not((layer0_outputs(783)) or (layer0_outputs(840)));
    outputs(2267) <= not((layer0_outputs(563)) xor (layer0_outputs(2526)));
    outputs(2268) <= (layer0_outputs(280)) and not (layer0_outputs(746));
    outputs(2269) <= layer0_outputs(1895);
    outputs(2270) <= (layer0_outputs(1115)) and (layer0_outputs(424));
    outputs(2271) <= layer0_outputs(2256);
    outputs(2272) <= (layer0_outputs(1284)) and not (layer0_outputs(1975));
    outputs(2273) <= (layer0_outputs(2279)) and not (layer0_outputs(1729));
    outputs(2274) <= (layer0_outputs(250)) and not (layer0_outputs(1898));
    outputs(2275) <= not((layer0_outputs(655)) or (layer0_outputs(3)));
    outputs(2276) <= not((layer0_outputs(72)) and (layer0_outputs(2144)));
    outputs(2277) <= not(layer0_outputs(1298));
    outputs(2278) <= not(layer0_outputs(541));
    outputs(2279) <= not(layer0_outputs(2240)) or (layer0_outputs(1021));
    outputs(2280) <= (layer0_outputs(964)) xor (layer0_outputs(1737));
    outputs(2281) <= (layer0_outputs(2521)) or (layer0_outputs(1192));
    outputs(2282) <= not(layer0_outputs(2458));
    outputs(2283) <= layer0_outputs(446);
    outputs(2284) <= (layer0_outputs(1979)) and (layer0_outputs(839));
    outputs(2285) <= not(layer0_outputs(75));
    outputs(2286) <= not(layer0_outputs(1360));
    outputs(2287) <= (layer0_outputs(2299)) and not (layer0_outputs(2074));
    outputs(2288) <= layer0_outputs(944);
    outputs(2289) <= not(layer0_outputs(359));
    outputs(2290) <= not(layer0_outputs(1852)) or (layer0_outputs(2501));
    outputs(2291) <= not((layer0_outputs(2493)) and (layer0_outputs(1631)));
    outputs(2292) <= not((layer0_outputs(1721)) xor (layer0_outputs(1012)));
    outputs(2293) <= not(layer0_outputs(113));
    outputs(2294) <= layer0_outputs(785);
    outputs(2295) <= layer0_outputs(258);
    outputs(2296) <= not((layer0_outputs(2197)) xor (layer0_outputs(1373)));
    outputs(2297) <= not(layer0_outputs(841));
    outputs(2298) <= not((layer0_outputs(45)) and (layer0_outputs(1216)));
    outputs(2299) <= (layer0_outputs(2489)) and not (layer0_outputs(2392));
    outputs(2300) <= (layer0_outputs(224)) and (layer0_outputs(1930));
    outputs(2301) <= layer0_outputs(2060);
    outputs(2302) <= layer0_outputs(63);
    outputs(2303) <= layer0_outputs(561);
    outputs(2304) <= layer0_outputs(2495);
    outputs(2305) <= (layer0_outputs(368)) and not (layer0_outputs(1817));
    outputs(2306) <= not(layer0_outputs(1378));
    outputs(2307) <= not((layer0_outputs(1085)) xor (layer0_outputs(1725)));
    outputs(2308) <= (layer0_outputs(1225)) and not (layer0_outputs(120));
    outputs(2309) <= not(layer0_outputs(1891));
    outputs(2310) <= not(layer0_outputs(948));
    outputs(2311) <= (layer0_outputs(204)) and not (layer0_outputs(830));
    outputs(2312) <= (layer0_outputs(177)) or (layer0_outputs(855));
    outputs(2313) <= not(layer0_outputs(2508));
    outputs(2314) <= (layer0_outputs(1915)) and not (layer0_outputs(2053));
    outputs(2315) <= (layer0_outputs(2363)) xor (layer0_outputs(2498));
    outputs(2316) <= not((layer0_outputs(1517)) xor (layer0_outputs(336)));
    outputs(2317) <= (layer0_outputs(363)) and not (layer0_outputs(1970));
    outputs(2318) <= layer0_outputs(462);
    outputs(2319) <= layer0_outputs(104);
    outputs(2320) <= not(layer0_outputs(502)) or (layer0_outputs(2055));
    outputs(2321) <= not((layer0_outputs(810)) or (layer0_outputs(1864)));
    outputs(2322) <= not((layer0_outputs(109)) xor (layer0_outputs(855)));
    outputs(2323) <= (layer0_outputs(1281)) and not (layer0_outputs(1030));
    outputs(2324) <= (layer0_outputs(1648)) xor (layer0_outputs(1867));
    outputs(2325) <= (layer0_outputs(2189)) xor (layer0_outputs(2450));
    outputs(2326) <= not((layer0_outputs(1705)) xor (layer0_outputs(1592)));
    outputs(2327) <= not(layer0_outputs(2547));
    outputs(2328) <= layer0_outputs(150);
    outputs(2329) <= layer0_outputs(2039);
    outputs(2330) <= not((layer0_outputs(761)) or (layer0_outputs(2440)));
    outputs(2331) <= layer0_outputs(2186);
    outputs(2332) <= layer0_outputs(599);
    outputs(2333) <= not(layer0_outputs(843)) or (layer0_outputs(544));
    outputs(2334) <= not(layer0_outputs(1633)) or (layer0_outputs(492));
    outputs(2335) <= layer0_outputs(1840);
    outputs(2336) <= not(layer0_outputs(1457));
    outputs(2337) <= (layer0_outputs(1735)) and not (layer0_outputs(1386));
    outputs(2338) <= (layer0_outputs(1250)) and (layer0_outputs(1742));
    outputs(2339) <= layer0_outputs(1662);
    outputs(2340) <= (layer0_outputs(1680)) xor (layer0_outputs(1857));
    outputs(2341) <= not(layer0_outputs(2447));
    outputs(2342) <= (layer0_outputs(503)) and not (layer0_outputs(1219));
    outputs(2343) <= (layer0_outputs(1685)) and not (layer0_outputs(2479));
    outputs(2344) <= (layer0_outputs(1889)) and not (layer0_outputs(2459));
    outputs(2345) <= not(layer0_outputs(2375)) or (layer0_outputs(672));
    outputs(2346) <= not(layer0_outputs(1068));
    outputs(2347) <= not(layer0_outputs(356));
    outputs(2348) <= layer0_outputs(743);
    outputs(2349) <= not(layer0_outputs(298));
    outputs(2350) <= not((layer0_outputs(505)) xor (layer0_outputs(1939)));
    outputs(2351) <= (layer0_outputs(3)) and not (layer0_outputs(2201));
    outputs(2352) <= (layer0_outputs(16)) and not (layer0_outputs(470));
    outputs(2353) <= (layer0_outputs(1109)) xor (layer0_outputs(135));
    outputs(2354) <= (layer0_outputs(1999)) and not (layer0_outputs(495));
    outputs(2355) <= (layer0_outputs(1890)) xor (layer0_outputs(851));
    outputs(2356) <= (layer0_outputs(425)) and not (layer0_outputs(1677));
    outputs(2357) <= not((layer0_outputs(1065)) xor (layer0_outputs(1338)));
    outputs(2358) <= not(layer0_outputs(1066));
    outputs(2359) <= (layer0_outputs(38)) and not (layer0_outputs(1637));
    outputs(2360) <= (layer0_outputs(1085)) and not (layer0_outputs(1308));
    outputs(2361) <= not(layer0_outputs(1348));
    outputs(2362) <= not(layer0_outputs(1386));
    outputs(2363) <= not(layer0_outputs(1434));
    outputs(2364) <= not((layer0_outputs(2471)) xor (layer0_outputs(127)));
    outputs(2365) <= layer0_outputs(2367);
    outputs(2366) <= layer0_outputs(2417);
    outputs(2367) <= layer0_outputs(2291);
    outputs(2368) <= (layer0_outputs(2555)) or (layer0_outputs(396));
    outputs(2369) <= (layer0_outputs(66)) and not (layer0_outputs(1194));
    outputs(2370) <= (layer0_outputs(750)) and not (layer0_outputs(2361));
    outputs(2371) <= not(layer0_outputs(52)) or (layer0_outputs(2357));
    outputs(2372) <= layer0_outputs(454);
    outputs(2373) <= (layer0_outputs(2136)) and not (layer0_outputs(1420));
    outputs(2374) <= not(layer0_outputs(729));
    outputs(2375) <= (layer0_outputs(2000)) xor (layer0_outputs(1994));
    outputs(2376) <= (layer0_outputs(892)) and (layer0_outputs(2149));
    outputs(2377) <= not(layer0_outputs(1815));
    outputs(2378) <= not(layer0_outputs(2031));
    outputs(2379) <= (layer0_outputs(1462)) and not (layer0_outputs(2316));
    outputs(2380) <= not((layer0_outputs(1447)) or (layer0_outputs(1532)));
    outputs(2381) <= layer0_outputs(1376);
    outputs(2382) <= (layer0_outputs(2077)) and not (layer0_outputs(2094));
    outputs(2383) <= not(layer0_outputs(215));
    outputs(2384) <= (layer0_outputs(2302)) and (layer0_outputs(484));
    outputs(2385) <= not(layer0_outputs(1382));
    outputs(2386) <= not(layer0_outputs(1343));
    outputs(2387) <= (layer0_outputs(1485)) and not (layer0_outputs(622));
    outputs(2388) <= (layer0_outputs(1965)) xor (layer0_outputs(2437));
    outputs(2389) <= not(layer0_outputs(2122));
    outputs(2390) <= layer0_outputs(707);
    outputs(2391) <= not(layer0_outputs(984));
    outputs(2392) <= not(layer0_outputs(2298));
    outputs(2393) <= layer0_outputs(651);
    outputs(2394) <= (layer0_outputs(2370)) and not (layer0_outputs(1768));
    outputs(2395) <= (layer0_outputs(1101)) and not (layer0_outputs(207));
    outputs(2396) <= not(layer0_outputs(2322));
    outputs(2397) <= not(layer0_outputs(1769));
    outputs(2398) <= (layer0_outputs(2388)) and not (layer0_outputs(227));
    outputs(2399) <= (layer0_outputs(1094)) xor (layer0_outputs(2509));
    outputs(2400) <= layer0_outputs(676);
    outputs(2401) <= (layer0_outputs(1667)) and (layer0_outputs(849));
    outputs(2402) <= (layer0_outputs(1602)) or (layer0_outputs(691));
    outputs(2403) <= (layer0_outputs(2378)) and (layer0_outputs(1013));
    outputs(2404) <= not(layer0_outputs(1658)) or (layer0_outputs(938));
    outputs(2405) <= not(layer0_outputs(1274));
    outputs(2406) <= (layer0_outputs(1842)) and not (layer0_outputs(2461));
    outputs(2407) <= not(layer0_outputs(1282));
    outputs(2408) <= not(layer0_outputs(1417)) or (layer0_outputs(1952));
    outputs(2409) <= (layer0_outputs(907)) or (layer0_outputs(723));
    outputs(2410) <= not((layer0_outputs(1757)) or (layer0_outputs(256)));
    outputs(2411) <= not(layer0_outputs(2007)) or (layer0_outputs(2387));
    outputs(2412) <= layer0_outputs(1698);
    outputs(2413) <= not(layer0_outputs(746)) or (layer0_outputs(598));
    outputs(2414) <= not(layer0_outputs(2391));
    outputs(2415) <= not((layer0_outputs(703)) or (layer0_outputs(2168)));
    outputs(2416) <= (layer0_outputs(2488)) and not (layer0_outputs(2227));
    outputs(2417) <= (layer0_outputs(2265)) and (layer0_outputs(1510));
    outputs(2418) <= not(layer0_outputs(434));
    outputs(2419) <= (layer0_outputs(902)) xor (layer0_outputs(1832));
    outputs(2420) <= not((layer0_outputs(380)) and (layer0_outputs(1469)));
    outputs(2421) <= (layer0_outputs(1534)) and not (layer0_outputs(1049));
    outputs(2422) <= not((layer0_outputs(1152)) or (layer0_outputs(1637)));
    outputs(2423) <= (layer0_outputs(895)) xor (layer0_outputs(2233));
    outputs(2424) <= (layer0_outputs(123)) and not (layer0_outputs(335));
    outputs(2425) <= not(layer0_outputs(261));
    outputs(2426) <= (layer0_outputs(2147)) and not (layer0_outputs(467));
    outputs(2427) <= (layer0_outputs(748)) and not (layer0_outputs(2050));
    outputs(2428) <= not((layer0_outputs(2468)) xor (layer0_outputs(1174)));
    outputs(2429) <= (layer0_outputs(724)) and (layer0_outputs(2202));
    outputs(2430) <= not(layer0_outputs(1317));
    outputs(2431) <= not(layer0_outputs(898));
    outputs(2432) <= not(layer0_outputs(87)) or (layer0_outputs(1238));
    outputs(2433) <= (layer0_outputs(1574)) and not (layer0_outputs(604));
    outputs(2434) <= (layer0_outputs(775)) or (layer0_outputs(1125));
    outputs(2435) <= layer0_outputs(1498);
    outputs(2436) <= not(layer0_outputs(1535));
    outputs(2437) <= not((layer0_outputs(1833)) or (layer0_outputs(1237)));
    outputs(2438) <= not(layer0_outputs(2326));
    outputs(2439) <= layer0_outputs(1442);
    outputs(2440) <= layer0_outputs(93);
    outputs(2441) <= not(layer0_outputs(2281));
    outputs(2442) <= not((layer0_outputs(0)) xor (layer0_outputs(1968)));
    outputs(2443) <= (layer0_outputs(302)) and not (layer0_outputs(342));
    outputs(2444) <= (layer0_outputs(1339)) xor (layer0_outputs(961));
    outputs(2445) <= (layer0_outputs(1357)) and (layer0_outputs(568));
    outputs(2446) <= not(layer0_outputs(2013));
    outputs(2447) <= (layer0_outputs(2519)) and not (layer0_outputs(1605));
    outputs(2448) <= (layer0_outputs(1143)) and not (layer0_outputs(2138));
    outputs(2449) <= not((layer0_outputs(755)) or (layer0_outputs(2252)));
    outputs(2450) <= not((layer0_outputs(2027)) xor (layer0_outputs(1007)));
    outputs(2451) <= (layer0_outputs(70)) and (layer0_outputs(1634));
    outputs(2452) <= not(layer0_outputs(33));
    outputs(2453) <= (layer0_outputs(90)) and (layer0_outputs(79));
    outputs(2454) <= layer0_outputs(291);
    outputs(2455) <= (layer0_outputs(1767)) or (layer0_outputs(1167));
    outputs(2456) <= not((layer0_outputs(336)) xor (layer0_outputs(124)));
    outputs(2457) <= (layer0_outputs(1790)) and (layer0_outputs(219));
    outputs(2458) <= (layer0_outputs(2525)) and (layer0_outputs(2274));
    outputs(2459) <= not((layer0_outputs(795)) or (layer0_outputs(2358)));
    outputs(2460) <= (layer0_outputs(250)) and (layer0_outputs(2551));
    outputs(2461) <= not(layer0_outputs(1982));
    outputs(2462) <= (layer0_outputs(1477)) and not (layer0_outputs(1444));
    outputs(2463) <= (layer0_outputs(2402)) and not (layer0_outputs(920));
    outputs(2464) <= (layer0_outputs(373)) and not (layer0_outputs(1252));
    outputs(2465) <= (layer0_outputs(15)) and not (layer0_outputs(2166));
    outputs(2466) <= not(layer0_outputs(489));
    outputs(2467) <= (layer0_outputs(2449)) and (layer0_outputs(2198));
    outputs(2468) <= not(layer0_outputs(22));
    outputs(2469) <= layer0_outputs(980);
    outputs(2470) <= (layer0_outputs(2499)) and not (layer0_outputs(2287));
    outputs(2471) <= layer0_outputs(105);
    outputs(2472) <= (layer0_outputs(2171)) and (layer0_outputs(2443));
    outputs(2473) <= (layer0_outputs(923)) and not (layer0_outputs(1064));
    outputs(2474) <= not((layer0_outputs(68)) and (layer0_outputs(2550)));
    outputs(2475) <= (layer0_outputs(762)) and not (layer0_outputs(2366));
    outputs(2476) <= (layer0_outputs(1937)) and (layer0_outputs(165));
    outputs(2477) <= (layer0_outputs(637)) xor (layer0_outputs(1256));
    outputs(2478) <= (layer0_outputs(799)) xor (layer0_outputs(1825));
    outputs(2479) <= not(layer0_outputs(1877)) or (layer0_outputs(499));
    outputs(2480) <= layer0_outputs(1325);
    outputs(2481) <= layer0_outputs(274);
    outputs(2482) <= layer0_outputs(1837);
    outputs(2483) <= layer0_outputs(2008);
    outputs(2484) <= (layer0_outputs(1423)) xor (layer0_outputs(1587));
    outputs(2485) <= not(layer0_outputs(1004));
    outputs(2486) <= not(layer0_outputs(2036));
    outputs(2487) <= not((layer0_outputs(1359)) or (layer0_outputs(2531)));
    outputs(2488) <= not(layer0_outputs(1150));
    outputs(2489) <= layer0_outputs(2169);
    outputs(2490) <= not(layer0_outputs(1035));
    outputs(2491) <= '1';
    outputs(2492) <= (layer0_outputs(2394)) and not (layer0_outputs(1128));
    outputs(2493) <= (layer0_outputs(628)) or (layer0_outputs(44));
    outputs(2494) <= (layer0_outputs(1990)) and not (layer0_outputs(30));
    outputs(2495) <= (layer0_outputs(653)) and not (layer0_outputs(481));
    outputs(2496) <= not(layer0_outputs(67));
    outputs(2497) <= not(layer0_outputs(767));
    outputs(2498) <= (layer0_outputs(1663)) and (layer0_outputs(2064));
    outputs(2499) <= (layer0_outputs(1490)) and not (layer0_outputs(2333));
    outputs(2500) <= not(layer0_outputs(1385));
    outputs(2501) <= not(layer0_outputs(547)) or (layer0_outputs(829));
    outputs(2502) <= not(layer0_outputs(2447)) or (layer0_outputs(1088));
    outputs(2503) <= not((layer0_outputs(1730)) or (layer0_outputs(2435)));
    outputs(2504) <= not(layer0_outputs(1812)) or (layer0_outputs(561));
    outputs(2505) <= not(layer0_outputs(1982));
    outputs(2506) <= layer0_outputs(2089);
    outputs(2507) <= not(layer0_outputs(261));
    outputs(2508) <= layer0_outputs(1957);
    outputs(2509) <= (layer0_outputs(1813)) and (layer0_outputs(533));
    outputs(2510) <= layer0_outputs(2311);
    outputs(2511) <= (layer0_outputs(192)) and not (layer0_outputs(471));
    outputs(2512) <= (layer0_outputs(294)) xor (layer0_outputs(2132));
    outputs(2513) <= not((layer0_outputs(218)) or (layer0_outputs(2385)));
    outputs(2514) <= (layer0_outputs(1582)) and not (layer0_outputs(1800));
    outputs(2515) <= not((layer0_outputs(2199)) xor (layer0_outputs(1278)));
    outputs(2516) <= layer0_outputs(907);
    outputs(2517) <= layer0_outputs(278);
    outputs(2518) <= not((layer0_outputs(2175)) or (layer0_outputs(1211)));
    outputs(2519) <= (layer0_outputs(2473)) and not (layer0_outputs(56));
    outputs(2520) <= layer0_outputs(1154);
    outputs(2521) <= not((layer0_outputs(725)) xor (layer0_outputs(554)));
    outputs(2522) <= (layer0_outputs(1540)) and (layer0_outputs(1731));
    outputs(2523) <= layer0_outputs(2346);
    outputs(2524) <= (layer0_outputs(2011)) and not (layer0_outputs(2466));
    outputs(2525) <= (layer0_outputs(1147)) or (layer0_outputs(2365));
    outputs(2526) <= not((layer0_outputs(1317)) or (layer0_outputs(1481)));
    outputs(2527) <= not((layer0_outputs(1952)) or (layer0_outputs(1261)));
    outputs(2528) <= not((layer0_outputs(1455)) or (layer0_outputs(704)));
    outputs(2529) <= (layer0_outputs(184)) and (layer0_outputs(1213));
    outputs(2530) <= not(layer0_outputs(825)) or (layer0_outputs(1405));
    outputs(2531) <= not(layer0_outputs(1736));
    outputs(2532) <= (layer0_outputs(682)) xor (layer0_outputs(2259));
    outputs(2533) <= not(layer0_outputs(74));
    outputs(2534) <= not(layer0_outputs(1434)) or (layer0_outputs(1613));
    outputs(2535) <= (layer0_outputs(1184)) and not (layer0_outputs(2251));
    outputs(2536) <= (layer0_outputs(331)) and not (layer0_outputs(449));
    outputs(2537) <= not(layer0_outputs(981));
    outputs(2538) <= not((layer0_outputs(804)) and (layer0_outputs(1735)));
    outputs(2539) <= (layer0_outputs(1556)) xor (layer0_outputs(603));
    outputs(2540) <= layer0_outputs(235);
    outputs(2541) <= not(layer0_outputs(1348));
    outputs(2542) <= layer0_outputs(100);
    outputs(2543) <= not((layer0_outputs(1968)) xor (layer0_outputs(2313)));
    outputs(2544) <= (layer0_outputs(486)) xor (layer0_outputs(32));
    outputs(2545) <= layer0_outputs(1170);
    outputs(2546) <= not(layer0_outputs(1792)) or (layer0_outputs(594));
    outputs(2547) <= (layer0_outputs(2146)) and not (layer0_outputs(253));
    outputs(2548) <= (layer0_outputs(1522)) and not (layer0_outputs(179));
    outputs(2549) <= not((layer0_outputs(2135)) or (layer0_outputs(1384)));
    outputs(2550) <= (layer0_outputs(636)) and (layer0_outputs(809));
    outputs(2551) <= not((layer0_outputs(39)) and (layer0_outputs(1535)));
    outputs(2552) <= not(layer0_outputs(577));
    outputs(2553) <= (layer0_outputs(1081)) and not (layer0_outputs(1423));
    outputs(2554) <= (layer0_outputs(1673)) and not (layer0_outputs(1885));
    outputs(2555) <= not((layer0_outputs(121)) or (layer0_outputs(2020)));
    outputs(2556) <= not(layer0_outputs(2007));
    outputs(2557) <= (layer0_outputs(1682)) and not (layer0_outputs(2191));
    outputs(2558) <= layer0_outputs(453);
    outputs(2559) <= layer0_outputs(2255);

end Behavioral;
