library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity logic_network is
    port (
        inputs : in std_logic_vector(255 downto 0);
        outputs : out std_logic_vector(10239 downto 0)
    );
end logic_network;

architecture Behavioral of logic_network is
    signal layer0_outputs : std_logic_vector(10239 downto 0);
    signal layer1_outputs : std_logic_vector(10239 downto 0);
    signal layer2_outputs : std_logic_vector(10239 downto 0);

begin

    layer0_outputs(0) <= (inputs(111)) and (inputs(75));
    layer0_outputs(1) <= (inputs(215)) or (inputs(254));
    layer0_outputs(2) <= (inputs(97)) and not (inputs(177));
    layer0_outputs(3) <= '1';
    layer0_outputs(4) <= (inputs(220)) and (inputs(216));
    layer0_outputs(5) <= not(inputs(164));
    layer0_outputs(6) <= inputs(95);
    layer0_outputs(7) <= inputs(72);
    layer0_outputs(8) <= inputs(181);
    layer0_outputs(9) <= not(inputs(109));
    layer0_outputs(10) <= not((inputs(37)) xor (inputs(19)));
    layer0_outputs(11) <= (inputs(250)) or (inputs(185));
    layer0_outputs(12) <= (inputs(48)) and not (inputs(124));
    layer0_outputs(13) <= '0';
    layer0_outputs(14) <= not((inputs(32)) or (inputs(201)));
    layer0_outputs(15) <= inputs(203);
    layer0_outputs(16) <= not((inputs(111)) or (inputs(51)));
    layer0_outputs(17) <= (inputs(46)) or (inputs(5));
    layer0_outputs(18) <= (inputs(34)) and not (inputs(59));
    layer0_outputs(19) <= inputs(87);
    layer0_outputs(20) <= inputs(199);
    layer0_outputs(21) <= '1';
    layer0_outputs(22) <= not(inputs(164));
    layer0_outputs(23) <= not(inputs(24)) or (inputs(182));
    layer0_outputs(24) <= not(inputs(245));
    layer0_outputs(25) <= inputs(227);
    layer0_outputs(26) <= not(inputs(40));
    layer0_outputs(27) <= not(inputs(183)) or (inputs(30));
    layer0_outputs(28) <= inputs(169);
    layer0_outputs(29) <= not(inputs(77));
    layer0_outputs(30) <= not((inputs(65)) or (inputs(151)));
    layer0_outputs(31) <= not(inputs(136));
    layer0_outputs(32) <= not(inputs(195)) or (inputs(71));
    layer0_outputs(33) <= (inputs(35)) or (inputs(44));
    layer0_outputs(34) <= (inputs(19)) and not (inputs(79));
    layer0_outputs(35) <= inputs(20);
    layer0_outputs(36) <= inputs(214);
    layer0_outputs(37) <= (inputs(35)) or (inputs(180));
    layer0_outputs(38) <= (inputs(249)) or (inputs(193));
    layer0_outputs(39) <= inputs(38);
    layer0_outputs(40) <= (inputs(138)) or (inputs(10));
    layer0_outputs(41) <= (inputs(105)) and not (inputs(240));
    layer0_outputs(42) <= inputs(91);
    layer0_outputs(43) <= inputs(213);
    layer0_outputs(44) <= (inputs(97)) or (inputs(107));
    layer0_outputs(45) <= not((inputs(111)) or (inputs(250)));
    layer0_outputs(46) <= not((inputs(174)) or (inputs(196)));
    layer0_outputs(47) <= not(inputs(183));
    layer0_outputs(48) <= inputs(163);
    layer0_outputs(49) <= not(inputs(80));
    layer0_outputs(50) <= not(inputs(233));
    layer0_outputs(51) <= (inputs(51)) and not (inputs(76));
    layer0_outputs(52) <= (inputs(51)) xor (inputs(84));
    layer0_outputs(53) <= inputs(235);
    layer0_outputs(54) <= (inputs(172)) and not (inputs(72));
    layer0_outputs(55) <= (inputs(179)) and not (inputs(191));
    layer0_outputs(56) <= inputs(5);
    layer0_outputs(57) <= '1';
    layer0_outputs(58) <= not(inputs(168)) or (inputs(188));
    layer0_outputs(59) <= (inputs(78)) or (inputs(54));
    layer0_outputs(60) <= not(inputs(44));
    layer0_outputs(61) <= not(inputs(175));
    layer0_outputs(62) <= inputs(27);
    layer0_outputs(63) <= not((inputs(140)) or (inputs(113)));
    layer0_outputs(64) <= not((inputs(24)) or (inputs(7)));
    layer0_outputs(65) <= '1';
    layer0_outputs(66) <= not((inputs(214)) or (inputs(186)));
    layer0_outputs(67) <= inputs(1);
    layer0_outputs(68) <= not(inputs(76));
    layer0_outputs(69) <= not(inputs(83));
    layer0_outputs(70) <= not(inputs(164));
    layer0_outputs(71) <= not((inputs(35)) or (inputs(183)));
    layer0_outputs(72) <= not(inputs(231)) or (inputs(112));
    layer0_outputs(73) <= '0';
    layer0_outputs(74) <= inputs(250);
    layer0_outputs(75) <= inputs(246);
    layer0_outputs(76) <= not((inputs(14)) or (inputs(33)));
    layer0_outputs(77) <= not(inputs(194));
    layer0_outputs(78) <= '1';
    layer0_outputs(79) <= not((inputs(194)) or (inputs(230)));
    layer0_outputs(80) <= (inputs(79)) xor (inputs(10));
    layer0_outputs(81) <= not(inputs(165)) or (inputs(71));
    layer0_outputs(82) <= not(inputs(56));
    layer0_outputs(83) <= inputs(91);
    layer0_outputs(84) <= inputs(210);
    layer0_outputs(85) <= not((inputs(44)) or (inputs(92)));
    layer0_outputs(86) <= inputs(125);
    layer0_outputs(87) <= (inputs(59)) and (inputs(12));
    layer0_outputs(88) <= not(inputs(22));
    layer0_outputs(89) <= inputs(214);
    layer0_outputs(90) <= (inputs(60)) or (inputs(126));
    layer0_outputs(91) <= inputs(238);
    layer0_outputs(92) <= (inputs(222)) xor (inputs(64));
    layer0_outputs(93) <= not(inputs(94));
    layer0_outputs(94) <= inputs(158);
    layer0_outputs(95) <= (inputs(216)) or (inputs(57));
    layer0_outputs(96) <= not(inputs(137));
    layer0_outputs(97) <= (inputs(193)) or (inputs(37));
    layer0_outputs(98) <= not(inputs(228)) or (inputs(94));
    layer0_outputs(99) <= not((inputs(78)) or (inputs(25)));
    layer0_outputs(100) <= not(inputs(109)) or (inputs(221));
    layer0_outputs(101) <= inputs(23);
    layer0_outputs(102) <= (inputs(64)) xor (inputs(66));
    layer0_outputs(103) <= (inputs(63)) xor (inputs(112));
    layer0_outputs(104) <= inputs(124);
    layer0_outputs(105) <= not(inputs(224)) or (inputs(193));
    layer0_outputs(106) <= '0';
    layer0_outputs(107) <= not((inputs(159)) or (inputs(23)));
    layer0_outputs(108) <= inputs(136);
    layer0_outputs(109) <= '1';
    layer0_outputs(110) <= (inputs(103)) and (inputs(44));
    layer0_outputs(111) <= '1';
    layer0_outputs(112) <= (inputs(22)) and (inputs(120));
    layer0_outputs(113) <= not(inputs(181)) or (inputs(35));
    layer0_outputs(114) <= '1';
    layer0_outputs(115) <= (inputs(167)) and (inputs(204));
    layer0_outputs(116) <= (inputs(91)) and not (inputs(112));
    layer0_outputs(117) <= (inputs(172)) xor (inputs(48));
    layer0_outputs(118) <= (inputs(249)) or (inputs(14));
    layer0_outputs(119) <= not((inputs(175)) or (inputs(233)));
    layer0_outputs(120) <= (inputs(33)) and not (inputs(137));
    layer0_outputs(121) <= not(inputs(4)) or (inputs(249));
    layer0_outputs(122) <= not(inputs(71));
    layer0_outputs(123) <= not(inputs(72));
    layer0_outputs(124) <= inputs(227);
    layer0_outputs(125) <= (inputs(157)) and not (inputs(208));
    layer0_outputs(126) <= not(inputs(19)) or (inputs(96));
    layer0_outputs(127) <= (inputs(70)) and not (inputs(146));
    layer0_outputs(128) <= not((inputs(204)) xor (inputs(228)));
    layer0_outputs(129) <= not(inputs(233));
    layer0_outputs(130) <= inputs(165);
    layer0_outputs(131) <= not(inputs(37));
    layer0_outputs(132) <= (inputs(49)) and (inputs(251));
    layer0_outputs(133) <= not((inputs(89)) xor (inputs(128)));
    layer0_outputs(134) <= not(inputs(231));
    layer0_outputs(135) <= (inputs(147)) xor (inputs(111));
    layer0_outputs(136) <= not((inputs(223)) or (inputs(163)));
    layer0_outputs(137) <= (inputs(43)) and (inputs(217));
    layer0_outputs(138) <= '1';
    layer0_outputs(139) <= (inputs(188)) and (inputs(90));
    layer0_outputs(140) <= inputs(179);
    layer0_outputs(141) <= inputs(208);
    layer0_outputs(142) <= (inputs(154)) and not (inputs(177));
    layer0_outputs(143) <= not((inputs(32)) and (inputs(102)));
    layer0_outputs(144) <= (inputs(151)) and not (inputs(129));
    layer0_outputs(145) <= (inputs(232)) xor (inputs(42));
    layer0_outputs(146) <= inputs(205);
    layer0_outputs(147) <= not((inputs(12)) or (inputs(50)));
    layer0_outputs(148) <= (inputs(149)) and not (inputs(15));
    layer0_outputs(149) <= not(inputs(229));
    layer0_outputs(150) <= (inputs(21)) and not (inputs(172));
    layer0_outputs(151) <= not((inputs(9)) and (inputs(72)));
    layer0_outputs(152) <= not(inputs(215)) or (inputs(100));
    layer0_outputs(153) <= (inputs(128)) and not (inputs(43));
    layer0_outputs(154) <= not((inputs(99)) and (inputs(29)));
    layer0_outputs(155) <= not((inputs(24)) and (inputs(152)));
    layer0_outputs(156) <= (inputs(35)) or (inputs(234));
    layer0_outputs(157) <= '1';
    layer0_outputs(158) <= (inputs(213)) or (inputs(204));
    layer0_outputs(159) <= not(inputs(136));
    layer0_outputs(160) <= not(inputs(204)) or (inputs(127));
    layer0_outputs(161) <= '0';
    layer0_outputs(162) <= '1';
    layer0_outputs(163) <= not(inputs(151)) or (inputs(100));
    layer0_outputs(164) <= not(inputs(203));
    layer0_outputs(165) <= inputs(247);
    layer0_outputs(166) <= not(inputs(69)) or (inputs(164));
    layer0_outputs(167) <= inputs(123);
    layer0_outputs(168) <= (inputs(250)) or (inputs(226));
    layer0_outputs(169) <= inputs(43);
    layer0_outputs(170) <= not(inputs(221)) or (inputs(117));
    layer0_outputs(171) <= inputs(168);
    layer0_outputs(172) <= not((inputs(61)) and (inputs(149)));
    layer0_outputs(173) <= not((inputs(83)) and (inputs(57)));
    layer0_outputs(174) <= inputs(22);
    layer0_outputs(175) <= not(inputs(247)) or (inputs(254));
    layer0_outputs(176) <= (inputs(11)) or (inputs(213));
    layer0_outputs(177) <= inputs(83);
    layer0_outputs(178) <= not(inputs(120)) or (inputs(83));
    layer0_outputs(179) <= (inputs(23)) and not (inputs(198));
    layer0_outputs(180) <= not(inputs(219));
    layer0_outputs(181) <= not(inputs(251));
    layer0_outputs(182) <= (inputs(71)) xor (inputs(37));
    layer0_outputs(183) <= inputs(250);
    layer0_outputs(184) <= (inputs(13)) and (inputs(175));
    layer0_outputs(185) <= not((inputs(48)) xor (inputs(118)));
    layer0_outputs(186) <= (inputs(204)) or (inputs(11));
    layer0_outputs(187) <= (inputs(123)) xor (inputs(170));
    layer0_outputs(188) <= not(inputs(248)) or (inputs(1));
    layer0_outputs(189) <= not(inputs(69)) or (inputs(162));
    layer0_outputs(190) <= (inputs(253)) or (inputs(47));
    layer0_outputs(191) <= inputs(87);
    layer0_outputs(192) <= (inputs(180)) or (inputs(61));
    layer0_outputs(193) <= not((inputs(24)) or (inputs(9)));
    layer0_outputs(194) <= not(inputs(252)) or (inputs(79));
    layer0_outputs(195) <= inputs(92);
    layer0_outputs(196) <= not(inputs(53)) or (inputs(141));
    layer0_outputs(197) <= inputs(43);
    layer0_outputs(198) <= not(inputs(179));
    layer0_outputs(199) <= not(inputs(212));
    layer0_outputs(200) <= (inputs(168)) and (inputs(88));
    layer0_outputs(201) <= (inputs(14)) xor (inputs(174));
    layer0_outputs(202) <= inputs(61);
    layer0_outputs(203) <= not(inputs(125));
    layer0_outputs(204) <= (inputs(101)) and not (inputs(48));
    layer0_outputs(205) <= (inputs(216)) and (inputs(110));
    layer0_outputs(206) <= not(inputs(175));
    layer0_outputs(207) <= not(inputs(45));
    layer0_outputs(208) <= not(inputs(98));
    layer0_outputs(209) <= (inputs(18)) or (inputs(140));
    layer0_outputs(210) <= not(inputs(36)) or (inputs(199));
    layer0_outputs(211) <= (inputs(42)) or (inputs(159));
    layer0_outputs(212) <= inputs(206);
    layer0_outputs(213) <= (inputs(83)) or (inputs(159));
    layer0_outputs(214) <= inputs(163);
    layer0_outputs(215) <= (inputs(103)) and not (inputs(97));
    layer0_outputs(216) <= not((inputs(122)) xor (inputs(223)));
    layer0_outputs(217) <= inputs(68);
    layer0_outputs(218) <= not(inputs(127));
    layer0_outputs(219) <= (inputs(165)) or (inputs(238));
    layer0_outputs(220) <= (inputs(213)) and not (inputs(61));
    layer0_outputs(221) <= not((inputs(42)) and (inputs(120)));
    layer0_outputs(222) <= not(inputs(51)) or (inputs(237));
    layer0_outputs(223) <= not((inputs(235)) or (inputs(86)));
    layer0_outputs(224) <= (inputs(145)) and not (inputs(167));
    layer0_outputs(225) <= not(inputs(88));
    layer0_outputs(226) <= '0';
    layer0_outputs(227) <= (inputs(29)) or (inputs(104));
    layer0_outputs(228) <= not(inputs(101));
    layer0_outputs(229) <= not(inputs(214)) or (inputs(30));
    layer0_outputs(230) <= inputs(162);
    layer0_outputs(231) <= not(inputs(106));
    layer0_outputs(232) <= (inputs(105)) and not (inputs(98));
    layer0_outputs(233) <= (inputs(181)) xor (inputs(204));
    layer0_outputs(234) <= not((inputs(9)) xor (inputs(33)));
    layer0_outputs(235) <= not(inputs(92)) or (inputs(1));
    layer0_outputs(236) <= not(inputs(82));
    layer0_outputs(237) <= not((inputs(5)) xor (inputs(157)));
    layer0_outputs(238) <= not(inputs(114));
    layer0_outputs(239) <= not(inputs(25));
    layer0_outputs(240) <= not(inputs(96));
    layer0_outputs(241) <= inputs(40);
    layer0_outputs(242) <= not((inputs(110)) xor (inputs(158)));
    layer0_outputs(243) <= inputs(219);
    layer0_outputs(244) <= '1';
    layer0_outputs(245) <= (inputs(177)) and not (inputs(112));
    layer0_outputs(246) <= '1';
    layer0_outputs(247) <= not((inputs(11)) or (inputs(179)));
    layer0_outputs(248) <= (inputs(3)) xor (inputs(237));
    layer0_outputs(249) <= not(inputs(197)) or (inputs(112));
    layer0_outputs(250) <= not((inputs(233)) or (inputs(234)));
    layer0_outputs(251) <= '1';
    layer0_outputs(252) <= not(inputs(92)) or (inputs(88));
    layer0_outputs(253) <= (inputs(82)) and not (inputs(235));
    layer0_outputs(254) <= (inputs(212)) or (inputs(238));
    layer0_outputs(255) <= (inputs(148)) and not (inputs(5));
    layer0_outputs(256) <= not(inputs(40)) or (inputs(129));
    layer0_outputs(257) <= (inputs(21)) and (inputs(188));
    layer0_outputs(258) <= not((inputs(94)) or (inputs(141)));
    layer0_outputs(259) <= inputs(76);
    layer0_outputs(260) <= (inputs(81)) and not (inputs(130));
    layer0_outputs(261) <= (inputs(168)) and not (inputs(249));
    layer0_outputs(262) <= not(inputs(212)) or (inputs(34));
    layer0_outputs(263) <= (inputs(153)) and not (inputs(198));
    layer0_outputs(264) <= inputs(191);
    layer0_outputs(265) <= not(inputs(58)) or (inputs(209));
    layer0_outputs(266) <= inputs(115);
    layer0_outputs(267) <= not(inputs(84));
    layer0_outputs(268) <= not(inputs(217)) or (inputs(139));
    layer0_outputs(269) <= not(inputs(247)) or (inputs(86));
    layer0_outputs(270) <= (inputs(112)) or (inputs(161));
    layer0_outputs(271) <= not((inputs(229)) or (inputs(146)));
    layer0_outputs(272) <= not(inputs(72));
    layer0_outputs(273) <= '1';
    layer0_outputs(274) <= not(inputs(77));
    layer0_outputs(275) <= inputs(90);
    layer0_outputs(276) <= inputs(162);
    layer0_outputs(277) <= not(inputs(173)) or (inputs(34));
    layer0_outputs(278) <= inputs(110);
    layer0_outputs(279) <= not((inputs(165)) or (inputs(101)));
    layer0_outputs(280) <= inputs(194);
    layer0_outputs(281) <= inputs(126);
    layer0_outputs(282) <= not(inputs(201)) or (inputs(122));
    layer0_outputs(283) <= not((inputs(195)) xor (inputs(168)));
    layer0_outputs(284) <= inputs(166);
    layer0_outputs(285) <= not(inputs(150));
    layer0_outputs(286) <= inputs(73);
    layer0_outputs(287) <= inputs(69);
    layer0_outputs(288) <= not(inputs(13));
    layer0_outputs(289) <= not(inputs(87)) or (inputs(34));
    layer0_outputs(290) <= not((inputs(186)) or (inputs(66)));
    layer0_outputs(291) <= inputs(201);
    layer0_outputs(292) <= not(inputs(245)) or (inputs(83));
    layer0_outputs(293) <= (inputs(184)) and not (inputs(9));
    layer0_outputs(294) <= (inputs(181)) xor (inputs(246));
    layer0_outputs(295) <= (inputs(39)) and not (inputs(180));
    layer0_outputs(296) <= (inputs(226)) or (inputs(32));
    layer0_outputs(297) <= (inputs(17)) or (inputs(32));
    layer0_outputs(298) <= not((inputs(166)) xor (inputs(89)));
    layer0_outputs(299) <= inputs(12);
    layer0_outputs(300) <= inputs(155);
    layer0_outputs(301) <= (inputs(32)) and not (inputs(29));
    layer0_outputs(302) <= inputs(169);
    layer0_outputs(303) <= not(inputs(132));
    layer0_outputs(304) <= not((inputs(125)) or (inputs(156)));
    layer0_outputs(305) <= not(inputs(178));
    layer0_outputs(306) <= not((inputs(28)) or (inputs(30)));
    layer0_outputs(307) <= not(inputs(56)) or (inputs(228));
    layer0_outputs(308) <= not(inputs(254)) or (inputs(57));
    layer0_outputs(309) <= inputs(182);
    layer0_outputs(310) <= not(inputs(119)) or (inputs(20));
    layer0_outputs(311) <= inputs(178);
    layer0_outputs(312) <= not(inputs(238));
    layer0_outputs(313) <= '0';
    layer0_outputs(314) <= (inputs(89)) and not (inputs(188));
    layer0_outputs(315) <= not(inputs(66)) or (inputs(16));
    layer0_outputs(316) <= (inputs(241)) and (inputs(223));
    layer0_outputs(317) <= not(inputs(25)) or (inputs(27));
    layer0_outputs(318) <= '1';
    layer0_outputs(319) <= (inputs(245)) and not (inputs(32));
    layer0_outputs(320) <= inputs(188);
    layer0_outputs(321) <= (inputs(226)) or (inputs(227));
    layer0_outputs(322) <= not((inputs(224)) or (inputs(56)));
    layer0_outputs(323) <= (inputs(44)) xor (inputs(76));
    layer0_outputs(324) <= (inputs(88)) or (inputs(10));
    layer0_outputs(325) <= not(inputs(62)) or (inputs(181));
    layer0_outputs(326) <= (inputs(173)) or (inputs(91));
    layer0_outputs(327) <= '0';
    layer0_outputs(328) <= not(inputs(215));
    layer0_outputs(329) <= (inputs(246)) and (inputs(220));
    layer0_outputs(330) <= not(inputs(241)) or (inputs(127));
    layer0_outputs(331) <= inputs(47);
    layer0_outputs(332) <= '0';
    layer0_outputs(333) <= not(inputs(66)) or (inputs(14));
    layer0_outputs(334) <= inputs(172);
    layer0_outputs(335) <= inputs(171);
    layer0_outputs(336) <= not(inputs(188));
    layer0_outputs(337) <= inputs(148);
    layer0_outputs(338) <= inputs(42);
    layer0_outputs(339) <= (inputs(147)) xor (inputs(85));
    layer0_outputs(340) <= not((inputs(100)) or (inputs(65)));
    layer0_outputs(341) <= (inputs(101)) and (inputs(164));
    layer0_outputs(342) <= inputs(169);
    layer0_outputs(343) <= not((inputs(69)) xor (inputs(219)));
    layer0_outputs(344) <= not((inputs(31)) and (inputs(210)));
    layer0_outputs(345) <= not(inputs(76)) or (inputs(202));
    layer0_outputs(346) <= inputs(77);
    layer0_outputs(347) <= (inputs(124)) or (inputs(53));
    layer0_outputs(348) <= (inputs(8)) or (inputs(45));
    layer0_outputs(349) <= '0';
    layer0_outputs(350) <= not(inputs(161)) or (inputs(88));
    layer0_outputs(351) <= not(inputs(105));
    layer0_outputs(352) <= not((inputs(88)) xor (inputs(161)));
    layer0_outputs(353) <= not((inputs(230)) xor (inputs(124)));
    layer0_outputs(354) <= not(inputs(56));
    layer0_outputs(355) <= not(inputs(237));
    layer0_outputs(356) <= not((inputs(88)) or (inputs(7)));
    layer0_outputs(357) <= not(inputs(242)) or (inputs(131));
    layer0_outputs(358) <= (inputs(198)) and not (inputs(178));
    layer0_outputs(359) <= not(inputs(1));
    layer0_outputs(360) <= not((inputs(193)) and (inputs(99)));
    layer0_outputs(361) <= inputs(114);
    layer0_outputs(362) <= not(inputs(58));
    layer0_outputs(363) <= not(inputs(133));
    layer0_outputs(364) <= (inputs(254)) or (inputs(63));
    layer0_outputs(365) <= (inputs(97)) xor (inputs(85));
    layer0_outputs(366) <= not(inputs(209));
    layer0_outputs(367) <= not((inputs(110)) and (inputs(244)));
    layer0_outputs(368) <= (inputs(63)) and not (inputs(33));
    layer0_outputs(369) <= (inputs(174)) xor (inputs(69));
    layer0_outputs(370) <= inputs(255);
    layer0_outputs(371) <= not(inputs(206));
    layer0_outputs(372) <= (inputs(36)) or (inputs(46));
    layer0_outputs(373) <= not(inputs(36));
    layer0_outputs(374) <= '0';
    layer0_outputs(375) <= (inputs(24)) or (inputs(27));
    layer0_outputs(376) <= inputs(178);
    layer0_outputs(377) <= not((inputs(97)) or (inputs(232)));
    layer0_outputs(378) <= not((inputs(227)) or (inputs(41)));
    layer0_outputs(379) <= inputs(94);
    layer0_outputs(380) <= not(inputs(240));
    layer0_outputs(381) <= (inputs(60)) or (inputs(189));
    layer0_outputs(382) <= not((inputs(46)) xor (inputs(227)));
    layer0_outputs(383) <= inputs(248);
    layer0_outputs(384) <= inputs(195);
    layer0_outputs(385) <= inputs(151);
    layer0_outputs(386) <= (inputs(151)) and not (inputs(193));
    layer0_outputs(387) <= inputs(214);
    layer0_outputs(388) <= (inputs(12)) xor (inputs(82));
    layer0_outputs(389) <= not((inputs(124)) or (inputs(75)));
    layer0_outputs(390) <= not((inputs(162)) or (inputs(163)));
    layer0_outputs(391) <= not((inputs(130)) or (inputs(154)));
    layer0_outputs(392) <= inputs(135);
    layer0_outputs(393) <= not(inputs(232));
    layer0_outputs(394) <= (inputs(218)) and not (inputs(27));
    layer0_outputs(395) <= not(inputs(109));
    layer0_outputs(396) <= not(inputs(184)) or (inputs(143));
    layer0_outputs(397) <= '1';
    layer0_outputs(398) <= not((inputs(180)) xor (inputs(206)));
    layer0_outputs(399) <= inputs(233);
    layer0_outputs(400) <= '0';
    layer0_outputs(401) <= (inputs(247)) or (inputs(58));
    layer0_outputs(402) <= (inputs(217)) and not (inputs(136));
    layer0_outputs(403) <= not((inputs(42)) or (inputs(226)));
    layer0_outputs(404) <= not(inputs(92)) or (inputs(79));
    layer0_outputs(405) <= not(inputs(158)) or (inputs(122));
    layer0_outputs(406) <= not(inputs(253));
    layer0_outputs(407) <= not(inputs(105));
    layer0_outputs(408) <= not((inputs(86)) xor (inputs(127)));
    layer0_outputs(409) <= not(inputs(16));
    layer0_outputs(410) <= not(inputs(108)) or (inputs(177));
    layer0_outputs(411) <= (inputs(231)) or (inputs(174));
    layer0_outputs(412) <= not(inputs(186)) or (inputs(30));
    layer0_outputs(413) <= inputs(75);
    layer0_outputs(414) <= (inputs(138)) and not (inputs(110));
    layer0_outputs(415) <= inputs(63);
    layer0_outputs(416) <= not(inputs(28)) or (inputs(220));
    layer0_outputs(417) <= not((inputs(49)) or (inputs(134)));
    layer0_outputs(418) <= not(inputs(71)) or (inputs(114));
    layer0_outputs(419) <= not((inputs(101)) or (inputs(178)));
    layer0_outputs(420) <= not(inputs(17));
    layer0_outputs(421) <= (inputs(83)) and (inputs(204));
    layer0_outputs(422) <= not((inputs(121)) or (inputs(180)));
    layer0_outputs(423) <= not((inputs(48)) and (inputs(48)));
    layer0_outputs(424) <= not(inputs(108));
    layer0_outputs(425) <= not(inputs(27)) or (inputs(223));
    layer0_outputs(426) <= not(inputs(0));
    layer0_outputs(427) <= not(inputs(17));
    layer0_outputs(428) <= not(inputs(233));
    layer0_outputs(429) <= inputs(132);
    layer0_outputs(430) <= not((inputs(43)) or (inputs(136)));
    layer0_outputs(431) <= inputs(23);
    layer0_outputs(432) <= not(inputs(170)) or (inputs(129));
    layer0_outputs(433) <= not(inputs(218)) or (inputs(68));
    layer0_outputs(434) <= (inputs(0)) and not (inputs(38));
    layer0_outputs(435) <= (inputs(94)) or (inputs(208));
    layer0_outputs(436) <= (inputs(204)) or (inputs(177));
    layer0_outputs(437) <= not(inputs(212));
    layer0_outputs(438) <= not((inputs(89)) and (inputs(7)));
    layer0_outputs(439) <= not(inputs(55));
    layer0_outputs(440) <= '1';
    layer0_outputs(441) <= inputs(103);
    layer0_outputs(442) <= (inputs(4)) xor (inputs(135));
    layer0_outputs(443) <= not((inputs(109)) xor (inputs(29)));
    layer0_outputs(444) <= not(inputs(161));
    layer0_outputs(445) <= (inputs(239)) or (inputs(131));
    layer0_outputs(446) <= not(inputs(99)) or (inputs(141));
    layer0_outputs(447) <= not((inputs(211)) xor (inputs(240)));
    layer0_outputs(448) <= not((inputs(239)) xor (inputs(170)));
    layer0_outputs(449) <= not((inputs(178)) or (inputs(168)));
    layer0_outputs(450) <= not((inputs(45)) or (inputs(97)));
    layer0_outputs(451) <= not(inputs(113));
    layer0_outputs(452) <= inputs(212);
    layer0_outputs(453) <= not((inputs(143)) or (inputs(180)));
    layer0_outputs(454) <= (inputs(113)) or (inputs(149));
    layer0_outputs(455) <= not(inputs(86));
    layer0_outputs(456) <= not(inputs(153));
    layer0_outputs(457) <= (inputs(52)) or (inputs(12));
    layer0_outputs(458) <= (inputs(48)) and not (inputs(42));
    layer0_outputs(459) <= inputs(57);
    layer0_outputs(460) <= not(inputs(35));
    layer0_outputs(461) <= (inputs(155)) and (inputs(44));
    layer0_outputs(462) <= inputs(228);
    layer0_outputs(463) <= inputs(248);
    layer0_outputs(464) <= not(inputs(7));
    layer0_outputs(465) <= (inputs(240)) and (inputs(170));
    layer0_outputs(466) <= not(inputs(106)) or (inputs(113));
    layer0_outputs(467) <= not(inputs(202)) or (inputs(94));
    layer0_outputs(468) <= not(inputs(59)) or (inputs(197));
    layer0_outputs(469) <= not((inputs(251)) xor (inputs(255)));
    layer0_outputs(470) <= not((inputs(24)) or (inputs(51)));
    layer0_outputs(471) <= inputs(229);
    layer0_outputs(472) <= inputs(232);
    layer0_outputs(473) <= not(inputs(149));
    layer0_outputs(474) <= (inputs(219)) or (inputs(255));
    layer0_outputs(475) <= (inputs(232)) and not (inputs(251));
    layer0_outputs(476) <= not(inputs(14));
    layer0_outputs(477) <= (inputs(172)) or (inputs(120));
    layer0_outputs(478) <= not(inputs(216)) or (inputs(229));
    layer0_outputs(479) <= (inputs(21)) or (inputs(124));
    layer0_outputs(480) <= not(inputs(117)) or (inputs(125));
    layer0_outputs(481) <= not((inputs(122)) or (inputs(40)));
    layer0_outputs(482) <= not(inputs(214));
    layer0_outputs(483) <= inputs(27);
    layer0_outputs(484) <= not((inputs(236)) and (inputs(144)));
    layer0_outputs(485) <= not(inputs(64)) or (inputs(56));
    layer0_outputs(486) <= inputs(141);
    layer0_outputs(487) <= (inputs(118)) and not (inputs(174));
    layer0_outputs(488) <= (inputs(43)) or (inputs(242));
    layer0_outputs(489) <= not((inputs(221)) xor (inputs(125)));
    layer0_outputs(490) <= not(inputs(247)) or (inputs(14));
    layer0_outputs(491) <= not(inputs(91));
    layer0_outputs(492) <= not(inputs(76));
    layer0_outputs(493) <= inputs(139);
    layer0_outputs(494) <= not(inputs(92));
    layer0_outputs(495) <= not((inputs(214)) or (inputs(106)));
    layer0_outputs(496) <= (inputs(202)) or (inputs(233));
    layer0_outputs(497) <= not(inputs(223));
    layer0_outputs(498) <= not((inputs(227)) or (inputs(211)));
    layer0_outputs(499) <= '0';
    layer0_outputs(500) <= inputs(49);
    layer0_outputs(501) <= not((inputs(110)) and (inputs(50)));
    layer0_outputs(502) <= not(inputs(137));
    layer0_outputs(503) <= not((inputs(147)) and (inputs(156)));
    layer0_outputs(504) <= (inputs(182)) or (inputs(127));
    layer0_outputs(505) <= inputs(247);
    layer0_outputs(506) <= (inputs(60)) and (inputs(97));
    layer0_outputs(507) <= not((inputs(48)) and (inputs(159)));
    layer0_outputs(508) <= not(inputs(53));
    layer0_outputs(509) <= not((inputs(2)) and (inputs(78)));
    layer0_outputs(510) <= (inputs(2)) and (inputs(186));
    layer0_outputs(511) <= (inputs(160)) or (inputs(143));
    layer0_outputs(512) <= (inputs(244)) and (inputs(246));
    layer0_outputs(513) <= inputs(210);
    layer0_outputs(514) <= (inputs(152)) and not (inputs(174));
    layer0_outputs(515) <= (inputs(63)) and not (inputs(99));
    layer0_outputs(516) <= (inputs(71)) and not (inputs(31));
    layer0_outputs(517) <= not(inputs(31));
    layer0_outputs(518) <= inputs(83);
    layer0_outputs(519) <= (inputs(79)) or (inputs(43));
    layer0_outputs(520) <= not(inputs(109)) or (inputs(252));
    layer0_outputs(521) <= inputs(119);
    layer0_outputs(522) <= (inputs(44)) and not (inputs(227));
    layer0_outputs(523) <= (inputs(255)) or (inputs(47));
    layer0_outputs(524) <= inputs(127);
    layer0_outputs(525) <= not(inputs(78)) or (inputs(15));
    layer0_outputs(526) <= (inputs(68)) and (inputs(61));
    layer0_outputs(527) <= not(inputs(15));
    layer0_outputs(528) <= (inputs(104)) xor (inputs(124));
    layer0_outputs(529) <= '1';
    layer0_outputs(530) <= (inputs(147)) or (inputs(173));
    layer0_outputs(531) <= (inputs(32)) xor (inputs(25));
    layer0_outputs(532) <= (inputs(180)) and not (inputs(45));
    layer0_outputs(533) <= inputs(84);
    layer0_outputs(534) <= (inputs(20)) and not (inputs(149));
    layer0_outputs(535) <= not((inputs(47)) or (inputs(115)));
    layer0_outputs(536) <= inputs(200);
    layer0_outputs(537) <= (inputs(48)) or (inputs(255));
    layer0_outputs(538) <= not(inputs(50)) or (inputs(74));
    layer0_outputs(539) <= (inputs(144)) xor (inputs(100));
    layer0_outputs(540) <= inputs(140);
    layer0_outputs(541) <= not(inputs(209));
    layer0_outputs(542) <= inputs(178);
    layer0_outputs(543) <= not((inputs(161)) xor (inputs(110)));
    layer0_outputs(544) <= not((inputs(82)) or (inputs(151)));
    layer0_outputs(545) <= (inputs(104)) and not (inputs(217));
    layer0_outputs(546) <= (inputs(145)) xor (inputs(13));
    layer0_outputs(547) <= inputs(12);
    layer0_outputs(548) <= (inputs(31)) and not (inputs(46));
    layer0_outputs(549) <= not(inputs(74));
    layer0_outputs(550) <= not((inputs(211)) or (inputs(142)));
    layer0_outputs(551) <= not(inputs(136)) or (inputs(64));
    layer0_outputs(552) <= not((inputs(49)) or (inputs(65)));
    layer0_outputs(553) <= not(inputs(2)) or (inputs(43));
    layer0_outputs(554) <= not(inputs(83));
    layer0_outputs(555) <= not((inputs(21)) xor (inputs(64)));
    layer0_outputs(556) <= not((inputs(17)) or (inputs(176)));
    layer0_outputs(557) <= not((inputs(210)) xor (inputs(102)));
    layer0_outputs(558) <= not(inputs(167)) or (inputs(43));
    layer0_outputs(559) <= not(inputs(13));
    layer0_outputs(560) <= inputs(83);
    layer0_outputs(561) <= not((inputs(223)) or (inputs(111)));
    layer0_outputs(562) <= not(inputs(32));
    layer0_outputs(563) <= inputs(30);
    layer0_outputs(564) <= not(inputs(101));
    layer0_outputs(565) <= inputs(217);
    layer0_outputs(566) <= not((inputs(52)) or (inputs(237)));
    layer0_outputs(567) <= not(inputs(127));
    layer0_outputs(568) <= not((inputs(223)) or (inputs(175)));
    layer0_outputs(569) <= not(inputs(162)) or (inputs(94));
    layer0_outputs(570) <= not(inputs(136));
    layer0_outputs(571) <= (inputs(119)) and not (inputs(49));
    layer0_outputs(572) <= '0';
    layer0_outputs(573) <= not((inputs(248)) xor (inputs(238)));
    layer0_outputs(574) <= not((inputs(89)) xor (inputs(117)));
    layer0_outputs(575) <= '0';
    layer0_outputs(576) <= (inputs(4)) xor (inputs(36));
    layer0_outputs(577) <= not(inputs(127));
    layer0_outputs(578) <= inputs(98);
    layer0_outputs(579) <= (inputs(67)) and not (inputs(74));
    layer0_outputs(580) <= inputs(87);
    layer0_outputs(581) <= not((inputs(154)) and (inputs(0)));
    layer0_outputs(582) <= (inputs(53)) and not (inputs(175));
    layer0_outputs(583) <= not((inputs(109)) xor (inputs(122)));
    layer0_outputs(584) <= not(inputs(114));
    layer0_outputs(585) <= not((inputs(210)) xor (inputs(148)));
    layer0_outputs(586) <= not((inputs(141)) or (inputs(8)));
    layer0_outputs(587) <= inputs(209);
    layer0_outputs(588) <= not(inputs(154)) or (inputs(227));
    layer0_outputs(589) <= (inputs(69)) and (inputs(153));
    layer0_outputs(590) <= not((inputs(70)) xor (inputs(67)));
    layer0_outputs(591) <= not(inputs(168));
    layer0_outputs(592) <= not((inputs(38)) xor (inputs(145)));
    layer0_outputs(593) <= '1';
    layer0_outputs(594) <= (inputs(161)) or (inputs(95));
    layer0_outputs(595) <= not((inputs(193)) xor (inputs(239)));
    layer0_outputs(596) <= inputs(89);
    layer0_outputs(597) <= inputs(33);
    layer0_outputs(598) <= not(inputs(141));
    layer0_outputs(599) <= (inputs(231)) or (inputs(65));
    layer0_outputs(600) <= not(inputs(119)) or (inputs(63));
    layer0_outputs(601) <= inputs(36);
    layer0_outputs(602) <= not((inputs(67)) xor (inputs(187)));
    layer0_outputs(603) <= not(inputs(240));
    layer0_outputs(604) <= not((inputs(126)) xor (inputs(109)));
    layer0_outputs(605) <= not((inputs(124)) or (inputs(35)));
    layer0_outputs(606) <= not((inputs(160)) or (inputs(239)));
    layer0_outputs(607) <= (inputs(166)) and not (inputs(129));
    layer0_outputs(608) <= '1';
    layer0_outputs(609) <= (inputs(107)) or (inputs(92));
    layer0_outputs(610) <= not(inputs(195));
    layer0_outputs(611) <= not(inputs(6)) or (inputs(68));
    layer0_outputs(612) <= not(inputs(64)) or (inputs(71));
    layer0_outputs(613) <= not((inputs(51)) or (inputs(123)));
    layer0_outputs(614) <= (inputs(100)) or (inputs(101));
    layer0_outputs(615) <= inputs(182);
    layer0_outputs(616) <= '0';
    layer0_outputs(617) <= not(inputs(20));
    layer0_outputs(618) <= not((inputs(9)) xor (inputs(15)));
    layer0_outputs(619) <= inputs(246);
    layer0_outputs(620) <= inputs(54);
    layer0_outputs(621) <= (inputs(125)) or (inputs(212));
    layer0_outputs(622) <= not((inputs(173)) or (inputs(207)));
    layer0_outputs(623) <= (inputs(56)) and not (inputs(240));
    layer0_outputs(624) <= not((inputs(198)) or (inputs(7)));
    layer0_outputs(625) <= inputs(233);
    layer0_outputs(626) <= inputs(126);
    layer0_outputs(627) <= inputs(77);
    layer0_outputs(628) <= not((inputs(225)) xor (inputs(216)));
    layer0_outputs(629) <= (inputs(171)) and not (inputs(62));
    layer0_outputs(630) <= not(inputs(6));
    layer0_outputs(631) <= '0';
    layer0_outputs(632) <= not(inputs(127));
    layer0_outputs(633) <= not((inputs(231)) and (inputs(61)));
    layer0_outputs(634) <= (inputs(141)) xor (inputs(176));
    layer0_outputs(635) <= not(inputs(213));
    layer0_outputs(636) <= not(inputs(158));
    layer0_outputs(637) <= not(inputs(116)) or (inputs(127));
    layer0_outputs(638) <= not(inputs(18));
    layer0_outputs(639) <= inputs(230);
    layer0_outputs(640) <= not(inputs(246));
    layer0_outputs(641) <= (inputs(1)) xor (inputs(24));
    layer0_outputs(642) <= (inputs(194)) and (inputs(141));
    layer0_outputs(643) <= (inputs(196)) and not (inputs(22));
    layer0_outputs(644) <= (inputs(59)) and not (inputs(140));
    layer0_outputs(645) <= (inputs(76)) and not (inputs(110));
    layer0_outputs(646) <= (inputs(203)) and not (inputs(229));
    layer0_outputs(647) <= '1';
    layer0_outputs(648) <= not((inputs(229)) and (inputs(158)));
    layer0_outputs(649) <= not(inputs(88));
    layer0_outputs(650) <= inputs(44);
    layer0_outputs(651) <= not((inputs(63)) xor (inputs(226)));
    layer0_outputs(652) <= (inputs(54)) and not (inputs(251));
    layer0_outputs(653) <= (inputs(254)) and not (inputs(232));
    layer0_outputs(654) <= not(inputs(151));
    layer0_outputs(655) <= (inputs(76)) xor (inputs(207));
    layer0_outputs(656) <= not((inputs(195)) xor (inputs(201)));
    layer0_outputs(657) <= not((inputs(172)) and (inputs(168)));
    layer0_outputs(658) <= '1';
    layer0_outputs(659) <= not(inputs(246)) or (inputs(146));
    layer0_outputs(660) <= inputs(168);
    layer0_outputs(661) <= not(inputs(234));
    layer0_outputs(662) <= not((inputs(64)) or (inputs(178)));
    layer0_outputs(663) <= (inputs(23)) or (inputs(195));
    layer0_outputs(664) <= not(inputs(212));
    layer0_outputs(665) <= not(inputs(118)) or (inputs(61));
    layer0_outputs(666) <= not(inputs(209)) or (inputs(138));
    layer0_outputs(667) <= (inputs(155)) and not (inputs(53));
    layer0_outputs(668) <= not((inputs(79)) xor (inputs(206)));
    layer0_outputs(669) <= (inputs(4)) and (inputs(130));
    layer0_outputs(670) <= inputs(11);
    layer0_outputs(671) <= not(inputs(252));
    layer0_outputs(672) <= not((inputs(212)) or (inputs(208)));
    layer0_outputs(673) <= (inputs(181)) and (inputs(176));
    layer0_outputs(674) <= not(inputs(122)) or (inputs(190));
    layer0_outputs(675) <= not((inputs(51)) or (inputs(14)));
    layer0_outputs(676) <= (inputs(214)) xor (inputs(81));
    layer0_outputs(677) <= not((inputs(211)) or (inputs(51)));
    layer0_outputs(678) <= not((inputs(209)) or (inputs(200)));
    layer0_outputs(679) <= (inputs(224)) or (inputs(94));
    layer0_outputs(680) <= not(inputs(173)) or (inputs(48));
    layer0_outputs(681) <= inputs(108);
    layer0_outputs(682) <= (inputs(125)) xor (inputs(233));
    layer0_outputs(683) <= not((inputs(11)) xor (inputs(127)));
    layer0_outputs(684) <= (inputs(150)) and not (inputs(123));
    layer0_outputs(685) <= not(inputs(186));
    layer0_outputs(686) <= (inputs(255)) xor (inputs(3));
    layer0_outputs(687) <= (inputs(108)) xor (inputs(18));
    layer0_outputs(688) <= not(inputs(78)) or (inputs(108));
    layer0_outputs(689) <= not(inputs(197));
    layer0_outputs(690) <= not(inputs(151));
    layer0_outputs(691) <= not(inputs(135)) or (inputs(141));
    layer0_outputs(692) <= inputs(139);
    layer0_outputs(693) <= not((inputs(29)) or (inputs(251)));
    layer0_outputs(694) <= not(inputs(135));
    layer0_outputs(695) <= inputs(5);
    layer0_outputs(696) <= (inputs(107)) and not (inputs(41));
    layer0_outputs(697) <= not((inputs(30)) or (inputs(7)));
    layer0_outputs(698) <= not((inputs(2)) or (inputs(66)));
    layer0_outputs(699) <= '0';
    layer0_outputs(700) <= not(inputs(17));
    layer0_outputs(701) <= (inputs(202)) or (inputs(60));
    layer0_outputs(702) <= inputs(96);
    layer0_outputs(703) <= (inputs(167)) and not (inputs(237));
    layer0_outputs(704) <= not(inputs(139)) or (inputs(9));
    layer0_outputs(705) <= (inputs(56)) and not (inputs(26));
    layer0_outputs(706) <= not(inputs(118));
    layer0_outputs(707) <= (inputs(27)) or (inputs(139));
    layer0_outputs(708) <= (inputs(94)) and (inputs(51));
    layer0_outputs(709) <= not(inputs(171));
    layer0_outputs(710) <= not(inputs(101));
    layer0_outputs(711) <= not(inputs(182)) or (inputs(10));
    layer0_outputs(712) <= (inputs(0)) xor (inputs(230));
    layer0_outputs(713) <= (inputs(198)) and not (inputs(171));
    layer0_outputs(714) <= not(inputs(85)) or (inputs(164));
    layer0_outputs(715) <= not((inputs(118)) xor (inputs(129)));
    layer0_outputs(716) <= not(inputs(74));
    layer0_outputs(717) <= not(inputs(163));
    layer0_outputs(718) <= not((inputs(245)) or (inputs(43)));
    layer0_outputs(719) <= not(inputs(248));
    layer0_outputs(720) <= inputs(83);
    layer0_outputs(721) <= (inputs(226)) or (inputs(34));
    layer0_outputs(722) <= '1';
    layer0_outputs(723) <= not((inputs(134)) xor (inputs(198)));
    layer0_outputs(724) <= (inputs(250)) and not (inputs(204));
    layer0_outputs(725) <= inputs(92);
    layer0_outputs(726) <= (inputs(66)) or (inputs(90));
    layer0_outputs(727) <= inputs(34);
    layer0_outputs(728) <= not(inputs(45)) or (inputs(27));
    layer0_outputs(729) <= (inputs(179)) and not (inputs(44));
    layer0_outputs(730) <= inputs(23);
    layer0_outputs(731) <= '1';
    layer0_outputs(732) <= inputs(158);
    layer0_outputs(733) <= not((inputs(192)) and (inputs(206)));
    layer0_outputs(734) <= (inputs(37)) and (inputs(52));
    layer0_outputs(735) <= '1';
    layer0_outputs(736) <= not((inputs(118)) xor (inputs(164)));
    layer0_outputs(737) <= (inputs(193)) or (inputs(68));
    layer0_outputs(738) <= (inputs(218)) or (inputs(128));
    layer0_outputs(739) <= '1';
    layer0_outputs(740) <= not((inputs(169)) or (inputs(3)));
    layer0_outputs(741) <= (inputs(112)) and not (inputs(255));
    layer0_outputs(742) <= not(inputs(81)) or (inputs(126));
    layer0_outputs(743) <= not((inputs(231)) or (inputs(116)));
    layer0_outputs(744) <= not((inputs(36)) or (inputs(18)));
    layer0_outputs(745) <= not(inputs(251)) or (inputs(236));
    layer0_outputs(746) <= not((inputs(211)) or (inputs(203)));
    layer0_outputs(747) <= inputs(246);
    layer0_outputs(748) <= not(inputs(116));
    layer0_outputs(749) <= not(inputs(208));
    layer0_outputs(750) <= not((inputs(226)) xor (inputs(211)));
    layer0_outputs(751) <= inputs(18);
    layer0_outputs(752) <= not(inputs(231));
    layer0_outputs(753) <= inputs(102);
    layer0_outputs(754) <= not(inputs(192));
    layer0_outputs(755) <= (inputs(19)) or (inputs(162));
    layer0_outputs(756) <= '0';
    layer0_outputs(757) <= (inputs(200)) and not (inputs(47));
    layer0_outputs(758) <= not((inputs(217)) xor (inputs(8)));
    layer0_outputs(759) <= not(inputs(132));
    layer0_outputs(760) <= not((inputs(79)) and (inputs(93)));
    layer0_outputs(761) <= (inputs(116)) or (inputs(141));
    layer0_outputs(762) <= inputs(182);
    layer0_outputs(763) <= '1';
    layer0_outputs(764) <= not(inputs(86)) or (inputs(107));
    layer0_outputs(765) <= not(inputs(139));
    layer0_outputs(766) <= inputs(60);
    layer0_outputs(767) <= inputs(148);
    layer0_outputs(768) <= not((inputs(230)) xor (inputs(247)));
    layer0_outputs(769) <= (inputs(53)) or (inputs(170));
    layer0_outputs(770) <= not((inputs(106)) xor (inputs(49)));
    layer0_outputs(771) <= (inputs(46)) xor (inputs(141));
    layer0_outputs(772) <= not(inputs(180));
    layer0_outputs(773) <= not(inputs(166));
    layer0_outputs(774) <= (inputs(76)) and not (inputs(189));
    layer0_outputs(775) <= (inputs(26)) and (inputs(203));
    layer0_outputs(776) <= '1';
    layer0_outputs(777) <= not(inputs(189)) or (inputs(195));
    layer0_outputs(778) <= not(inputs(163));
    layer0_outputs(779) <= not(inputs(27));
    layer0_outputs(780) <= not(inputs(22));
    layer0_outputs(781) <= (inputs(147)) or (inputs(38));
    layer0_outputs(782) <= not(inputs(7));
    layer0_outputs(783) <= not(inputs(126));
    layer0_outputs(784) <= not((inputs(57)) or (inputs(62)));
    layer0_outputs(785) <= inputs(135);
    layer0_outputs(786) <= not(inputs(122));
    layer0_outputs(787) <= (inputs(142)) and not (inputs(39));
    layer0_outputs(788) <= (inputs(230)) or (inputs(248));
    layer0_outputs(789) <= not(inputs(215)) or (inputs(49));
    layer0_outputs(790) <= not(inputs(180));
    layer0_outputs(791) <= not(inputs(241));
    layer0_outputs(792) <= (inputs(224)) and (inputs(139));
    layer0_outputs(793) <= (inputs(183)) or (inputs(148));
    layer0_outputs(794) <= not(inputs(81)) or (inputs(54));
    layer0_outputs(795) <= inputs(104);
    layer0_outputs(796) <= (inputs(155)) and not (inputs(223));
    layer0_outputs(797) <= (inputs(224)) or (inputs(133));
    layer0_outputs(798) <= inputs(204);
    layer0_outputs(799) <= not(inputs(103));
    layer0_outputs(800) <= not(inputs(42));
    layer0_outputs(801) <= inputs(11);
    layer0_outputs(802) <= '0';
    layer0_outputs(803) <= not((inputs(110)) or (inputs(93)));
    layer0_outputs(804) <= not(inputs(215));
    layer0_outputs(805) <= not(inputs(68));
    layer0_outputs(806) <= not(inputs(11));
    layer0_outputs(807) <= inputs(98);
    layer0_outputs(808) <= (inputs(6)) and not (inputs(29));
    layer0_outputs(809) <= (inputs(5)) and not (inputs(60));
    layer0_outputs(810) <= not(inputs(85));
    layer0_outputs(811) <= (inputs(22)) or (inputs(94));
    layer0_outputs(812) <= not((inputs(47)) xor (inputs(133)));
    layer0_outputs(813) <= (inputs(196)) or (inputs(10));
    layer0_outputs(814) <= (inputs(255)) or (inputs(95));
    layer0_outputs(815) <= not((inputs(223)) or (inputs(250)));
    layer0_outputs(816) <= not(inputs(28));
    layer0_outputs(817) <= (inputs(36)) and (inputs(67));
    layer0_outputs(818) <= not(inputs(184)) or (inputs(74));
    layer0_outputs(819) <= (inputs(25)) or (inputs(90));
    layer0_outputs(820) <= (inputs(243)) and not (inputs(6));
    layer0_outputs(821) <= (inputs(252)) or (inputs(164));
    layer0_outputs(822) <= (inputs(106)) xor (inputs(88));
    layer0_outputs(823) <= not(inputs(87));
    layer0_outputs(824) <= not(inputs(117));
    layer0_outputs(825) <= (inputs(102)) or (inputs(146));
    layer0_outputs(826) <= (inputs(222)) xor (inputs(127));
    layer0_outputs(827) <= (inputs(247)) and not (inputs(72));
    layer0_outputs(828) <= not(inputs(54)) or (inputs(124));
    layer0_outputs(829) <= '1';
    layer0_outputs(830) <= (inputs(119)) and (inputs(148));
    layer0_outputs(831) <= inputs(177);
    layer0_outputs(832) <= not(inputs(98)) or (inputs(192));
    layer0_outputs(833) <= inputs(152);
    layer0_outputs(834) <= not((inputs(68)) or (inputs(158)));
    layer0_outputs(835) <= (inputs(237)) and not (inputs(173));
    layer0_outputs(836) <= not((inputs(158)) and (inputs(41)));
    layer0_outputs(837) <= (inputs(83)) or (inputs(199));
    layer0_outputs(838) <= inputs(72);
    layer0_outputs(839) <= not(inputs(28));
    layer0_outputs(840) <= (inputs(233)) and not (inputs(248));
    layer0_outputs(841) <= inputs(152);
    layer0_outputs(842) <= (inputs(10)) and (inputs(116));
    layer0_outputs(843) <= not(inputs(10));
    layer0_outputs(844) <= (inputs(121)) or (inputs(82));
    layer0_outputs(845) <= (inputs(195)) or (inputs(62));
    layer0_outputs(846) <= inputs(105);
    layer0_outputs(847) <= (inputs(37)) or (inputs(6));
    layer0_outputs(848) <= (inputs(58)) xor (inputs(108));
    layer0_outputs(849) <= not(inputs(163));
    layer0_outputs(850) <= (inputs(116)) and (inputs(37));
    layer0_outputs(851) <= (inputs(17)) or (inputs(24));
    layer0_outputs(852) <= (inputs(170)) or (inputs(37));
    layer0_outputs(853) <= inputs(178);
    layer0_outputs(854) <= not(inputs(131)) or (inputs(34));
    layer0_outputs(855) <= not(inputs(21));
    layer0_outputs(856) <= '0';
    layer0_outputs(857) <= not((inputs(53)) and (inputs(39)));
    layer0_outputs(858) <= not((inputs(42)) xor (inputs(73)));
    layer0_outputs(859) <= not(inputs(56)) or (inputs(219));
    layer0_outputs(860) <= inputs(115);
    layer0_outputs(861) <= not((inputs(199)) or (inputs(245)));
    layer0_outputs(862) <= (inputs(110)) or (inputs(164));
    layer0_outputs(863) <= (inputs(195)) or (inputs(95));
    layer0_outputs(864) <= '1';
    layer0_outputs(865) <= '1';
    layer0_outputs(866) <= not(inputs(74)) or (inputs(111));
    layer0_outputs(867) <= (inputs(186)) and not (inputs(5));
    layer0_outputs(868) <= not(inputs(166));
    layer0_outputs(869) <= inputs(216);
    layer0_outputs(870) <= inputs(144);
    layer0_outputs(871) <= inputs(97);
    layer0_outputs(872) <= inputs(9);
    layer0_outputs(873) <= not((inputs(168)) or (inputs(32)));
    layer0_outputs(874) <= (inputs(223)) and not (inputs(250));
    layer0_outputs(875) <= not((inputs(238)) or (inputs(113)));
    layer0_outputs(876) <= not(inputs(220));
    layer0_outputs(877) <= (inputs(18)) and (inputs(171));
    layer0_outputs(878) <= not(inputs(154)) or (inputs(174));
    layer0_outputs(879) <= not(inputs(162)) or (inputs(192));
    layer0_outputs(880) <= not(inputs(102));
    layer0_outputs(881) <= not(inputs(175)) or (inputs(193));
    layer0_outputs(882) <= not(inputs(29));
    layer0_outputs(883) <= inputs(249);
    layer0_outputs(884) <= not(inputs(209)) or (inputs(224));
    layer0_outputs(885) <= inputs(231);
    layer0_outputs(886) <= not(inputs(10)) or (inputs(145));
    layer0_outputs(887) <= not(inputs(215));
    layer0_outputs(888) <= (inputs(113)) or (inputs(72));
    layer0_outputs(889) <= not(inputs(236));
    layer0_outputs(890) <= (inputs(184)) and not (inputs(225));
    layer0_outputs(891) <= not((inputs(196)) or (inputs(14)));
    layer0_outputs(892) <= (inputs(160)) or (inputs(207));
    layer0_outputs(893) <= '1';
    layer0_outputs(894) <= (inputs(177)) xor (inputs(0));
    layer0_outputs(895) <= (inputs(70)) and not (inputs(143));
    layer0_outputs(896) <= (inputs(23)) and (inputs(28));
    layer0_outputs(897) <= not(inputs(6)) or (inputs(98));
    layer0_outputs(898) <= '0';
    layer0_outputs(899) <= (inputs(120)) and not (inputs(14));
    layer0_outputs(900) <= inputs(222);
    layer0_outputs(901) <= not(inputs(215)) or (inputs(137));
    layer0_outputs(902) <= not(inputs(20));
    layer0_outputs(903) <= not(inputs(158)) or (inputs(41));
    layer0_outputs(904) <= not((inputs(248)) or (inputs(9)));
    layer0_outputs(905) <= (inputs(146)) and not (inputs(15));
    layer0_outputs(906) <= '0';
    layer0_outputs(907) <= not((inputs(68)) xor (inputs(80)));
    layer0_outputs(908) <= inputs(177);
    layer0_outputs(909) <= not((inputs(19)) and (inputs(107)));
    layer0_outputs(910) <= not((inputs(190)) xor (inputs(140)));
    layer0_outputs(911) <= not((inputs(11)) and (inputs(207)));
    layer0_outputs(912) <= not((inputs(154)) xor (inputs(241)));
    layer0_outputs(913) <= not(inputs(188)) or (inputs(55));
    layer0_outputs(914) <= (inputs(204)) and not (inputs(145));
    layer0_outputs(915) <= not(inputs(22));
    layer0_outputs(916) <= (inputs(203)) or (inputs(190));
    layer0_outputs(917) <= not(inputs(210));
    layer0_outputs(918) <= inputs(242);
    layer0_outputs(919) <= not(inputs(19)) or (inputs(175));
    layer0_outputs(920) <= not((inputs(97)) or (inputs(180)));
    layer0_outputs(921) <= (inputs(44)) and not (inputs(89));
    layer0_outputs(922) <= not(inputs(213));
    layer0_outputs(923) <= (inputs(250)) xor (inputs(24));
    layer0_outputs(924) <= (inputs(172)) xor (inputs(205));
    layer0_outputs(925) <= not(inputs(7)) or (inputs(247));
    layer0_outputs(926) <= inputs(210);
    layer0_outputs(927) <= not(inputs(209)) or (inputs(210));
    layer0_outputs(928) <= not(inputs(168));
    layer0_outputs(929) <= not(inputs(230));
    layer0_outputs(930) <= not((inputs(48)) or (inputs(120)));
    layer0_outputs(931) <= (inputs(49)) xor (inputs(94));
    layer0_outputs(932) <= not(inputs(68)) or (inputs(63));
    layer0_outputs(933) <= not(inputs(23)) or (inputs(16));
    layer0_outputs(934) <= (inputs(105)) and not (inputs(63));
    layer0_outputs(935) <= not(inputs(182));
    layer0_outputs(936) <= not((inputs(75)) and (inputs(156)));
    layer0_outputs(937) <= not((inputs(201)) or (inputs(130)));
    layer0_outputs(938) <= (inputs(204)) and (inputs(159));
    layer0_outputs(939) <= not((inputs(48)) or (inputs(199)));
    layer0_outputs(940) <= not((inputs(216)) or (inputs(177)));
    layer0_outputs(941) <= (inputs(140)) and (inputs(50));
    layer0_outputs(942) <= (inputs(53)) or (inputs(134));
    layer0_outputs(943) <= not((inputs(48)) or (inputs(66)));
    layer0_outputs(944) <= not(inputs(30));
    layer0_outputs(945) <= '1';
    layer0_outputs(946) <= (inputs(223)) and not (inputs(176));
    layer0_outputs(947) <= (inputs(57)) or (inputs(176));
    layer0_outputs(948) <= not(inputs(122)) or (inputs(249));
    layer0_outputs(949) <= inputs(220);
    layer0_outputs(950) <= inputs(153);
    layer0_outputs(951) <= (inputs(80)) or (inputs(150));
    layer0_outputs(952) <= not(inputs(97)) or (inputs(255));
    layer0_outputs(953) <= (inputs(153)) or (inputs(97));
    layer0_outputs(954) <= inputs(133);
    layer0_outputs(955) <= inputs(163);
    layer0_outputs(956) <= not(inputs(110));
    layer0_outputs(957) <= not(inputs(107));
    layer0_outputs(958) <= not((inputs(207)) or (inputs(174)));
    layer0_outputs(959) <= not((inputs(255)) or (inputs(51)));
    layer0_outputs(960) <= inputs(229);
    layer0_outputs(961) <= '1';
    layer0_outputs(962) <= inputs(164);
    layer0_outputs(963) <= (inputs(92)) xor (inputs(116));
    layer0_outputs(964) <= inputs(80);
    layer0_outputs(965) <= (inputs(184)) and not (inputs(81));
    layer0_outputs(966) <= not((inputs(180)) and (inputs(229)));
    layer0_outputs(967) <= not(inputs(51));
    layer0_outputs(968) <= not(inputs(31)) or (inputs(124));
    layer0_outputs(969) <= not((inputs(12)) and (inputs(46)));
    layer0_outputs(970) <= not(inputs(112)) or (inputs(176));
    layer0_outputs(971) <= not(inputs(122));
    layer0_outputs(972) <= (inputs(169)) or (inputs(47));
    layer0_outputs(973) <= inputs(230);
    layer0_outputs(974) <= not(inputs(37));
    layer0_outputs(975) <= not(inputs(155)) or (inputs(84));
    layer0_outputs(976) <= inputs(229);
    layer0_outputs(977) <= inputs(146);
    layer0_outputs(978) <= inputs(82);
    layer0_outputs(979) <= (inputs(172)) and not (inputs(107));
    layer0_outputs(980) <= not((inputs(82)) and (inputs(96)));
    layer0_outputs(981) <= not((inputs(118)) or (inputs(120)));
    layer0_outputs(982) <= (inputs(33)) xor (inputs(137));
    layer0_outputs(983) <= '1';
    layer0_outputs(984) <= not(inputs(32));
    layer0_outputs(985) <= not((inputs(58)) and (inputs(69)));
    layer0_outputs(986) <= (inputs(190)) and not (inputs(71));
    layer0_outputs(987) <= (inputs(118)) xor (inputs(196));
    layer0_outputs(988) <= (inputs(65)) xor (inputs(76));
    layer0_outputs(989) <= not((inputs(238)) or (inputs(101)));
    layer0_outputs(990) <= not((inputs(34)) or (inputs(64)));
    layer0_outputs(991) <= (inputs(15)) or (inputs(2));
    layer0_outputs(992) <= inputs(184);
    layer0_outputs(993) <= inputs(60);
    layer0_outputs(994) <= not((inputs(170)) or (inputs(90)));
    layer0_outputs(995) <= not((inputs(164)) and (inputs(58)));
    layer0_outputs(996) <= not(inputs(120)) or (inputs(206));
    layer0_outputs(997) <= (inputs(36)) or (inputs(32));
    layer0_outputs(998) <= not((inputs(235)) or (inputs(147)));
    layer0_outputs(999) <= not((inputs(72)) xor (inputs(43)));
    layer0_outputs(1000) <= not((inputs(115)) or (inputs(30)));
    layer0_outputs(1001) <= (inputs(26)) xor (inputs(224));
    layer0_outputs(1002) <= inputs(70);
    layer0_outputs(1003) <= not(inputs(12)) or (inputs(255));
    layer0_outputs(1004) <= (inputs(176)) and not (inputs(15));
    layer0_outputs(1005) <= (inputs(195)) and not (inputs(30));
    layer0_outputs(1006) <= (inputs(188)) or (inputs(228));
    layer0_outputs(1007) <= not(inputs(123)) or (inputs(201));
    layer0_outputs(1008) <= (inputs(13)) xor (inputs(177));
    layer0_outputs(1009) <= inputs(25);
    layer0_outputs(1010) <= not(inputs(102));
    layer0_outputs(1011) <= not((inputs(38)) or (inputs(126)));
    layer0_outputs(1012) <= not(inputs(95));
    layer0_outputs(1013) <= inputs(110);
    layer0_outputs(1014) <= inputs(22);
    layer0_outputs(1015) <= not((inputs(163)) or (inputs(150)));
    layer0_outputs(1016) <= (inputs(33)) or (inputs(14));
    layer0_outputs(1017) <= not(inputs(166));
    layer0_outputs(1018) <= inputs(129);
    layer0_outputs(1019) <= '1';
    layer0_outputs(1020) <= inputs(147);
    layer0_outputs(1021) <= (inputs(191)) and not (inputs(189));
    layer0_outputs(1022) <= not(inputs(215)) or (inputs(87));
    layer0_outputs(1023) <= (inputs(215)) or (inputs(128));
    layer0_outputs(1024) <= not(inputs(67));
    layer0_outputs(1025) <= inputs(70);
    layer0_outputs(1026) <= not(inputs(115));
    layer0_outputs(1027) <= (inputs(130)) xor (inputs(101));
    layer0_outputs(1028) <= (inputs(213)) and not (inputs(27));
    layer0_outputs(1029) <= not(inputs(211));
    layer0_outputs(1030) <= inputs(113);
    layer0_outputs(1031) <= not((inputs(69)) or (inputs(218)));
    layer0_outputs(1032) <= not(inputs(10)) or (inputs(14));
    layer0_outputs(1033) <= not((inputs(245)) xor (inputs(91)));
    layer0_outputs(1034) <= inputs(23);
    layer0_outputs(1035) <= (inputs(89)) and not (inputs(248));
    layer0_outputs(1036) <= not(inputs(169));
    layer0_outputs(1037) <= inputs(202);
    layer0_outputs(1038) <= (inputs(5)) and not (inputs(107));
    layer0_outputs(1039) <= (inputs(62)) xor (inputs(13));
    layer0_outputs(1040) <= inputs(9);
    layer0_outputs(1041) <= not((inputs(76)) and (inputs(68)));
    layer0_outputs(1042) <= (inputs(33)) or (inputs(157));
    layer0_outputs(1043) <= (inputs(18)) or (inputs(215));
    layer0_outputs(1044) <= (inputs(216)) or (inputs(246));
    layer0_outputs(1045) <= not(inputs(25)) or (inputs(52));
    layer0_outputs(1046) <= (inputs(39)) xor (inputs(142));
    layer0_outputs(1047) <= inputs(101);
    layer0_outputs(1048) <= not((inputs(92)) xor (inputs(27)));
    layer0_outputs(1049) <= not(inputs(183)) or (inputs(97));
    layer0_outputs(1050) <= (inputs(178)) and not (inputs(137));
    layer0_outputs(1051) <= not(inputs(255));
    layer0_outputs(1052) <= inputs(78);
    layer0_outputs(1053) <= (inputs(22)) or (inputs(6));
    layer0_outputs(1054) <= not((inputs(72)) xor (inputs(8)));
    layer0_outputs(1055) <= not(inputs(91)) or (inputs(69));
    layer0_outputs(1056) <= not((inputs(15)) or (inputs(138)));
    layer0_outputs(1057) <= inputs(171);
    layer0_outputs(1058) <= not((inputs(49)) xor (inputs(242)));
    layer0_outputs(1059) <= (inputs(173)) and not (inputs(2));
    layer0_outputs(1060) <= (inputs(94)) xor (inputs(211));
    layer0_outputs(1061) <= not((inputs(98)) xor (inputs(98)));
    layer0_outputs(1062) <= not(inputs(138));
    layer0_outputs(1063) <= not(inputs(53));
    layer0_outputs(1064) <= not(inputs(67)) or (inputs(201));
    layer0_outputs(1065) <= (inputs(201)) or (inputs(101));
    layer0_outputs(1066) <= inputs(145);
    layer0_outputs(1067) <= not(inputs(175));
    layer0_outputs(1068) <= (inputs(180)) and not (inputs(88));
    layer0_outputs(1069) <= (inputs(161)) and (inputs(70));
    layer0_outputs(1070) <= (inputs(201)) or (inputs(162));
    layer0_outputs(1071) <= (inputs(82)) and not (inputs(78));
    layer0_outputs(1072) <= (inputs(248)) or (inputs(142));
    layer0_outputs(1073) <= inputs(218);
    layer0_outputs(1074) <= inputs(8);
    layer0_outputs(1075) <= (inputs(164)) xor (inputs(160));
    layer0_outputs(1076) <= not(inputs(32)) or (inputs(57));
    layer0_outputs(1077) <= not(inputs(228)) or (inputs(175));
    layer0_outputs(1078) <= not((inputs(131)) or (inputs(127)));
    layer0_outputs(1079) <= not(inputs(102));
    layer0_outputs(1080) <= not((inputs(79)) and (inputs(249)));
    layer0_outputs(1081) <= not(inputs(26)) or (inputs(157));
    layer0_outputs(1082) <= not(inputs(245)) or (inputs(147));
    layer0_outputs(1083) <= inputs(215);
    layer0_outputs(1084) <= (inputs(212)) and not (inputs(141));
    layer0_outputs(1085) <= '0';
    layer0_outputs(1086) <= (inputs(252)) and not (inputs(72));
    layer0_outputs(1087) <= inputs(83);
    layer0_outputs(1088) <= not(inputs(249)) or (inputs(102));
    layer0_outputs(1089) <= (inputs(58)) and not (inputs(52));
    layer0_outputs(1090) <= not((inputs(65)) xor (inputs(7)));
    layer0_outputs(1091) <= (inputs(121)) or (inputs(65));
    layer0_outputs(1092) <= not(inputs(68)) or (inputs(32));
    layer0_outputs(1093) <= not(inputs(44));
    layer0_outputs(1094) <= (inputs(247)) and not (inputs(182));
    layer0_outputs(1095) <= not(inputs(60)) or (inputs(3));
    layer0_outputs(1096) <= inputs(75);
    layer0_outputs(1097) <= not(inputs(97));
    layer0_outputs(1098) <= inputs(216);
    layer0_outputs(1099) <= (inputs(243)) and not (inputs(156));
    layer0_outputs(1100) <= (inputs(125)) and not (inputs(211));
    layer0_outputs(1101) <= not((inputs(13)) xor (inputs(72)));
    layer0_outputs(1102) <= not((inputs(0)) or (inputs(95)));
    layer0_outputs(1103) <= (inputs(116)) or (inputs(153));
    layer0_outputs(1104) <= not(inputs(231));
    layer0_outputs(1105) <= not(inputs(26)) or (inputs(244));
    layer0_outputs(1106) <= (inputs(41)) or (inputs(94));
    layer0_outputs(1107) <= not((inputs(32)) or (inputs(194)));
    layer0_outputs(1108) <= inputs(208);
    layer0_outputs(1109) <= inputs(115);
    layer0_outputs(1110) <= (inputs(77)) and not (inputs(254));
    layer0_outputs(1111) <= (inputs(189)) and (inputs(51));
    layer0_outputs(1112) <= (inputs(183)) or (inputs(51));
    layer0_outputs(1113) <= (inputs(44)) and not (inputs(27));
    layer0_outputs(1114) <= (inputs(17)) or (inputs(74));
    layer0_outputs(1115) <= not(inputs(72));
    layer0_outputs(1116) <= inputs(230);
    layer0_outputs(1117) <= not(inputs(162));
    layer0_outputs(1118) <= not((inputs(189)) and (inputs(48)));
    layer0_outputs(1119) <= not((inputs(81)) or (inputs(116)));
    layer0_outputs(1120) <= inputs(104);
    layer0_outputs(1121) <= (inputs(160)) or (inputs(171));
    layer0_outputs(1122) <= inputs(234);
    layer0_outputs(1123) <= not(inputs(215));
    layer0_outputs(1124) <= (inputs(222)) and not (inputs(75));
    layer0_outputs(1125) <= not(inputs(101)) or (inputs(71));
    layer0_outputs(1126) <= not(inputs(117));
    layer0_outputs(1127) <= not(inputs(227)) or (inputs(213));
    layer0_outputs(1128) <= '0';
    layer0_outputs(1129) <= (inputs(56)) and (inputs(122));
    layer0_outputs(1130) <= not(inputs(15));
    layer0_outputs(1131) <= inputs(219);
    layer0_outputs(1132) <= not((inputs(197)) xor (inputs(42)));
    layer0_outputs(1133) <= not((inputs(23)) or (inputs(223)));
    layer0_outputs(1134) <= not(inputs(228));
    layer0_outputs(1135) <= inputs(36);
    layer0_outputs(1136) <= inputs(230);
    layer0_outputs(1137) <= inputs(189);
    layer0_outputs(1138) <= (inputs(141)) and (inputs(54));
    layer0_outputs(1139) <= (inputs(162)) xor (inputs(160));
    layer0_outputs(1140) <= not(inputs(64));
    layer0_outputs(1141) <= not((inputs(11)) and (inputs(65)));
    layer0_outputs(1142) <= (inputs(128)) and not (inputs(71));
    layer0_outputs(1143) <= (inputs(123)) or (inputs(51));
    layer0_outputs(1144) <= not((inputs(218)) or (inputs(202)));
    layer0_outputs(1145) <= inputs(1);
    layer0_outputs(1146) <= (inputs(116)) xor (inputs(1));
    layer0_outputs(1147) <= (inputs(136)) and not (inputs(226));
    layer0_outputs(1148) <= '0';
    layer0_outputs(1149) <= not(inputs(90));
    layer0_outputs(1150) <= not((inputs(204)) or (inputs(227)));
    layer0_outputs(1151) <= (inputs(122)) or (inputs(31));
    layer0_outputs(1152) <= (inputs(233)) and not (inputs(34));
    layer0_outputs(1153) <= not((inputs(143)) or (inputs(87)));
    layer0_outputs(1154) <= not((inputs(20)) or (inputs(209)));
    layer0_outputs(1155) <= (inputs(52)) or (inputs(40));
    layer0_outputs(1156) <= inputs(92);
    layer0_outputs(1157) <= not((inputs(19)) and (inputs(68)));
    layer0_outputs(1158) <= not((inputs(85)) xor (inputs(93)));
    layer0_outputs(1159) <= not(inputs(154)) or (inputs(9));
    layer0_outputs(1160) <= not((inputs(182)) xor (inputs(114)));
    layer0_outputs(1161) <= not((inputs(113)) or (inputs(134)));
    layer0_outputs(1162) <= (inputs(178)) and (inputs(163));
    layer0_outputs(1163) <= not((inputs(220)) xor (inputs(244)));
    layer0_outputs(1164) <= inputs(211);
    layer0_outputs(1165) <= not((inputs(185)) and (inputs(253)));
    layer0_outputs(1166) <= not(inputs(75));
    layer0_outputs(1167) <= inputs(68);
    layer0_outputs(1168) <= not(inputs(225)) or (inputs(112));
    layer0_outputs(1169) <= not(inputs(191));
    layer0_outputs(1170) <= not(inputs(87)) or (inputs(33));
    layer0_outputs(1171) <= not(inputs(29));
    layer0_outputs(1172) <= not((inputs(74)) or (inputs(94)));
    layer0_outputs(1173) <= not(inputs(126));
    layer0_outputs(1174) <= (inputs(154)) xor (inputs(42));
    layer0_outputs(1175) <= not(inputs(73));
    layer0_outputs(1176) <= '0';
    layer0_outputs(1177) <= not(inputs(78));
    layer0_outputs(1178) <= not(inputs(169)) or (inputs(98));
    layer0_outputs(1179) <= not(inputs(183));
    layer0_outputs(1180) <= not(inputs(76)) or (inputs(191));
    layer0_outputs(1181) <= not((inputs(61)) or (inputs(86)));
    layer0_outputs(1182) <= (inputs(200)) or (inputs(32));
    layer0_outputs(1183) <= (inputs(24)) and not (inputs(18));
    layer0_outputs(1184) <= (inputs(21)) and (inputs(14));
    layer0_outputs(1185) <= not((inputs(124)) and (inputs(223)));
    layer0_outputs(1186) <= (inputs(189)) or (inputs(46));
    layer0_outputs(1187) <= not(inputs(153));
    layer0_outputs(1188) <= inputs(82);
    layer0_outputs(1189) <= not((inputs(244)) and (inputs(97)));
    layer0_outputs(1190) <= '0';
    layer0_outputs(1191) <= not(inputs(90)) or (inputs(247));
    layer0_outputs(1192) <= not((inputs(188)) or (inputs(201)));
    layer0_outputs(1193) <= inputs(38);
    layer0_outputs(1194) <= inputs(71);
    layer0_outputs(1195) <= not(inputs(54));
    layer0_outputs(1196) <= not(inputs(33));
    layer0_outputs(1197) <= inputs(169);
    layer0_outputs(1198) <= (inputs(22)) or (inputs(121));
    layer0_outputs(1199) <= not((inputs(106)) or (inputs(114)));
    layer0_outputs(1200) <= not(inputs(180)) or (inputs(50));
    layer0_outputs(1201) <= not(inputs(230));
    layer0_outputs(1202) <= inputs(3);
    layer0_outputs(1203) <= inputs(128);
    layer0_outputs(1204) <= (inputs(97)) and not (inputs(69));
    layer0_outputs(1205) <= inputs(130);
    layer0_outputs(1206) <= (inputs(0)) xor (inputs(125));
    layer0_outputs(1207) <= (inputs(193)) xor (inputs(132));
    layer0_outputs(1208) <= not(inputs(156)) or (inputs(63));
    layer0_outputs(1209) <= (inputs(241)) and (inputs(64));
    layer0_outputs(1210) <= '0';
    layer0_outputs(1211) <= not(inputs(69)) or (inputs(147));
    layer0_outputs(1212) <= '0';
    layer0_outputs(1213) <= not(inputs(6));
    layer0_outputs(1214) <= (inputs(68)) or (inputs(101));
    layer0_outputs(1215) <= not(inputs(235));
    layer0_outputs(1216) <= not((inputs(174)) xor (inputs(208)));
    layer0_outputs(1217) <= inputs(180);
    layer0_outputs(1218) <= inputs(20);
    layer0_outputs(1219) <= not(inputs(193));
    layer0_outputs(1220) <= not(inputs(109)) or (inputs(235));
    layer0_outputs(1221) <= not(inputs(75));
    layer0_outputs(1222) <= (inputs(47)) or (inputs(80));
    layer0_outputs(1223) <= not((inputs(177)) or (inputs(141)));
    layer0_outputs(1224) <= not(inputs(71)) or (inputs(238));
    layer0_outputs(1225) <= inputs(121);
    layer0_outputs(1226) <= inputs(183);
    layer0_outputs(1227) <= inputs(246);
    layer0_outputs(1228) <= inputs(216);
    layer0_outputs(1229) <= (inputs(23)) and not (inputs(69));
    layer0_outputs(1230) <= (inputs(49)) and not (inputs(179));
    layer0_outputs(1231) <= not(inputs(98));
    layer0_outputs(1232) <= (inputs(219)) and not (inputs(67));
    layer0_outputs(1233) <= (inputs(169)) or (inputs(28));
    layer0_outputs(1234) <= not(inputs(221));
    layer0_outputs(1235) <= (inputs(198)) or (inputs(253));
    layer0_outputs(1236) <= not(inputs(228));
    layer0_outputs(1237) <= not(inputs(67)) or (inputs(217));
    layer0_outputs(1238) <= (inputs(132)) and not (inputs(212));
    layer0_outputs(1239) <= (inputs(45)) and not (inputs(86));
    layer0_outputs(1240) <= inputs(164);
    layer0_outputs(1241) <= (inputs(116)) and not (inputs(222));
    layer0_outputs(1242) <= not((inputs(175)) or (inputs(189)));
    layer0_outputs(1243) <= not(inputs(161));
    layer0_outputs(1244) <= (inputs(18)) and (inputs(221));
    layer0_outputs(1245) <= (inputs(40)) and (inputs(58));
    layer0_outputs(1246) <= (inputs(19)) or (inputs(187));
    layer0_outputs(1247) <= (inputs(81)) or (inputs(130));
    layer0_outputs(1248) <= not(inputs(155));
    layer0_outputs(1249) <= not(inputs(167));
    layer0_outputs(1250) <= (inputs(250)) and not (inputs(35));
    layer0_outputs(1251) <= not(inputs(58));
    layer0_outputs(1252) <= '1';
    layer0_outputs(1253) <= (inputs(232)) or (inputs(189));
    layer0_outputs(1254) <= not((inputs(182)) or (inputs(69)));
    layer0_outputs(1255) <= '1';
    layer0_outputs(1256) <= not((inputs(194)) or (inputs(216)));
    layer0_outputs(1257) <= inputs(52);
    layer0_outputs(1258) <= not((inputs(39)) or (inputs(197)));
    layer0_outputs(1259) <= (inputs(227)) and (inputs(146));
    layer0_outputs(1260) <= (inputs(78)) or (inputs(102));
    layer0_outputs(1261) <= not(inputs(122)) or (inputs(146));
    layer0_outputs(1262) <= inputs(102);
    layer0_outputs(1263) <= not((inputs(162)) or (inputs(171)));
    layer0_outputs(1264) <= (inputs(127)) xor (inputs(68));
    layer0_outputs(1265) <= inputs(176);
    layer0_outputs(1266) <= not(inputs(135)) or (inputs(216));
    layer0_outputs(1267) <= inputs(152);
    layer0_outputs(1268) <= (inputs(9)) and not (inputs(183));
    layer0_outputs(1269) <= inputs(101);
    layer0_outputs(1270) <= (inputs(206)) and not (inputs(145));
    layer0_outputs(1271) <= (inputs(91)) or (inputs(255));
    layer0_outputs(1272) <= (inputs(39)) xor (inputs(42));
    layer0_outputs(1273) <= inputs(135);
    layer0_outputs(1274) <= not((inputs(73)) or (inputs(187)));
    layer0_outputs(1275) <= not((inputs(232)) xor (inputs(126)));
    layer0_outputs(1276) <= not(inputs(211));
    layer0_outputs(1277) <= not((inputs(243)) and (inputs(106)));
    layer0_outputs(1278) <= inputs(150);
    layer0_outputs(1279) <= not((inputs(95)) xor (inputs(234)));
    layer0_outputs(1280) <= not(inputs(11)) or (inputs(170));
    layer0_outputs(1281) <= '1';
    layer0_outputs(1282) <= '1';
    layer0_outputs(1283) <= not((inputs(188)) xor (inputs(193)));
    layer0_outputs(1284) <= not(inputs(129));
    layer0_outputs(1285) <= inputs(70);
    layer0_outputs(1286) <= not(inputs(181)) or (inputs(247));
    layer0_outputs(1287) <= not((inputs(137)) or (inputs(109)));
    layer0_outputs(1288) <= not(inputs(248));
    layer0_outputs(1289) <= (inputs(155)) or (inputs(146));
    layer0_outputs(1290) <= not(inputs(22));
    layer0_outputs(1291) <= not(inputs(36)) or (inputs(85));
    layer0_outputs(1292) <= (inputs(111)) or (inputs(22));
    layer0_outputs(1293) <= not(inputs(80)) or (inputs(105));
    layer0_outputs(1294) <= (inputs(94)) xor (inputs(154));
    layer0_outputs(1295) <= inputs(173);
    layer0_outputs(1296) <= inputs(175);
    layer0_outputs(1297) <= not(inputs(228));
    layer0_outputs(1298) <= not((inputs(190)) or (inputs(61)));
    layer0_outputs(1299) <= not(inputs(110));
    layer0_outputs(1300) <= (inputs(219)) or (inputs(5));
    layer0_outputs(1301) <= not(inputs(180));
    layer0_outputs(1302) <= not(inputs(201)) or (inputs(30));
    layer0_outputs(1303) <= not((inputs(15)) xor (inputs(62)));
    layer0_outputs(1304) <= not((inputs(33)) or (inputs(107)));
    layer0_outputs(1305) <= not(inputs(78));
    layer0_outputs(1306) <= (inputs(85)) or (inputs(189));
    layer0_outputs(1307) <= inputs(70);
    layer0_outputs(1308) <= (inputs(64)) xor (inputs(34));
    layer0_outputs(1309) <= inputs(116);
    layer0_outputs(1310) <= not(inputs(179)) or (inputs(125));
    layer0_outputs(1311) <= not(inputs(136)) or (inputs(209));
    layer0_outputs(1312) <= (inputs(45)) xor (inputs(207));
    layer0_outputs(1313) <= (inputs(88)) and not (inputs(144));
    layer0_outputs(1314) <= '1';
    layer0_outputs(1315) <= not(inputs(250));
    layer0_outputs(1316) <= not((inputs(182)) or (inputs(108)));
    layer0_outputs(1317) <= (inputs(158)) xor (inputs(214));
    layer0_outputs(1318) <= inputs(87);
    layer0_outputs(1319) <= (inputs(189)) or (inputs(46));
    layer0_outputs(1320) <= inputs(78);
    layer0_outputs(1321) <= not(inputs(249));
    layer0_outputs(1322) <= not(inputs(99)) or (inputs(193));
    layer0_outputs(1323) <= inputs(98);
    layer0_outputs(1324) <= (inputs(9)) or (inputs(162));
    layer0_outputs(1325) <= not((inputs(5)) or (inputs(212)));
    layer0_outputs(1326) <= '1';
    layer0_outputs(1327) <= inputs(70);
    layer0_outputs(1328) <= (inputs(43)) xor (inputs(202));
    layer0_outputs(1329) <= (inputs(232)) xor (inputs(22));
    layer0_outputs(1330) <= inputs(41);
    layer0_outputs(1331) <= not(inputs(91));
    layer0_outputs(1332) <= not(inputs(10));
    layer0_outputs(1333) <= not((inputs(11)) xor (inputs(134)));
    layer0_outputs(1334) <= inputs(145);
    layer0_outputs(1335) <= inputs(249);
    layer0_outputs(1336) <= inputs(188);
    layer0_outputs(1337) <= (inputs(25)) or (inputs(54));
    layer0_outputs(1338) <= not((inputs(200)) xor (inputs(197)));
    layer0_outputs(1339) <= (inputs(215)) and not (inputs(99));
    layer0_outputs(1340) <= not((inputs(236)) xor (inputs(93)));
    layer0_outputs(1341) <= (inputs(219)) and not (inputs(143));
    layer0_outputs(1342) <= (inputs(213)) and not (inputs(73));
    layer0_outputs(1343) <= (inputs(251)) xor (inputs(148));
    layer0_outputs(1344) <= (inputs(132)) or (inputs(220));
    layer0_outputs(1345) <= (inputs(109)) and (inputs(120));
    layer0_outputs(1346) <= (inputs(176)) or (inputs(237));
    layer0_outputs(1347) <= inputs(165);
    layer0_outputs(1348) <= (inputs(189)) or (inputs(247));
    layer0_outputs(1349) <= not(inputs(230));
    layer0_outputs(1350) <= (inputs(95)) and not (inputs(74));
    layer0_outputs(1351) <= not((inputs(222)) or (inputs(190)));
    layer0_outputs(1352) <= not(inputs(59)) or (inputs(96));
    layer0_outputs(1353) <= not((inputs(76)) xor (inputs(3)));
    layer0_outputs(1354) <= (inputs(26)) and not (inputs(211));
    layer0_outputs(1355) <= not(inputs(147));
    layer0_outputs(1356) <= not((inputs(215)) xor (inputs(201)));
    layer0_outputs(1357) <= not(inputs(153));
    layer0_outputs(1358) <= (inputs(58)) or (inputs(43));
    layer0_outputs(1359) <= not(inputs(205)) or (inputs(18));
    layer0_outputs(1360) <= (inputs(250)) and not (inputs(138));
    layer0_outputs(1361) <= not(inputs(205)) or (inputs(32));
    layer0_outputs(1362) <= (inputs(40)) or (inputs(234));
    layer0_outputs(1363) <= not(inputs(183));
    layer0_outputs(1364) <= (inputs(38)) and not (inputs(51));
    layer0_outputs(1365) <= inputs(17);
    layer0_outputs(1366) <= (inputs(52)) and not (inputs(214));
    layer0_outputs(1367) <= inputs(153);
    layer0_outputs(1368) <= (inputs(227)) or (inputs(51));
    layer0_outputs(1369) <= (inputs(74)) and not (inputs(192));
    layer0_outputs(1370) <= not((inputs(199)) or (inputs(162)));
    layer0_outputs(1371) <= not((inputs(142)) or (inputs(141)));
    layer0_outputs(1372) <= inputs(150);
    layer0_outputs(1373) <= not((inputs(209)) or (inputs(199)));
    layer0_outputs(1374) <= (inputs(57)) and not (inputs(116));
    layer0_outputs(1375) <= not((inputs(161)) or (inputs(132)));
    layer0_outputs(1376) <= inputs(160);
    layer0_outputs(1377) <= '1';
    layer0_outputs(1378) <= not((inputs(57)) or (inputs(63)));
    layer0_outputs(1379) <= (inputs(172)) xor (inputs(104));
    layer0_outputs(1380) <= (inputs(71)) and not (inputs(46));
    layer0_outputs(1381) <= not(inputs(26)) or (inputs(191));
    layer0_outputs(1382) <= not(inputs(176));
    layer0_outputs(1383) <= (inputs(81)) and not (inputs(154));
    layer0_outputs(1384) <= inputs(214);
    layer0_outputs(1385) <= not(inputs(179));
    layer0_outputs(1386) <= not(inputs(165));
    layer0_outputs(1387) <= inputs(241);
    layer0_outputs(1388) <= not((inputs(37)) or (inputs(74)));
    layer0_outputs(1389) <= (inputs(148)) or (inputs(17));
    layer0_outputs(1390) <= '0';
    layer0_outputs(1391) <= not(inputs(194));
    layer0_outputs(1392) <= inputs(165);
    layer0_outputs(1393) <= not((inputs(184)) and (inputs(55)));
    layer0_outputs(1394) <= inputs(222);
    layer0_outputs(1395) <= not(inputs(77)) or (inputs(238));
    layer0_outputs(1396) <= not((inputs(32)) or (inputs(76)));
    layer0_outputs(1397) <= not(inputs(211));
    layer0_outputs(1398) <= (inputs(108)) and not (inputs(241));
    layer0_outputs(1399) <= not((inputs(98)) or (inputs(31)));
    layer0_outputs(1400) <= (inputs(129)) xor (inputs(161));
    layer0_outputs(1401) <= (inputs(38)) and not (inputs(204));
    layer0_outputs(1402) <= (inputs(166)) and (inputs(15));
    layer0_outputs(1403) <= (inputs(199)) and not (inputs(100));
    layer0_outputs(1404) <= not((inputs(37)) or (inputs(123)));
    layer0_outputs(1405) <= inputs(117);
    layer0_outputs(1406) <= inputs(115);
    layer0_outputs(1407) <= (inputs(74)) or (inputs(54));
    layer0_outputs(1408) <= (inputs(89)) and not (inputs(233));
    layer0_outputs(1409) <= inputs(41);
    layer0_outputs(1410) <= (inputs(78)) or (inputs(226));
    layer0_outputs(1411) <= '1';
    layer0_outputs(1412) <= not(inputs(181)) or (inputs(204));
    layer0_outputs(1413) <= (inputs(22)) and not (inputs(127));
    layer0_outputs(1414) <= (inputs(183)) xor (inputs(224));
    layer0_outputs(1415) <= not(inputs(132));
    layer0_outputs(1416) <= not(inputs(230));
    layer0_outputs(1417) <= not(inputs(39)) or (inputs(97));
    layer0_outputs(1418) <= (inputs(158)) xor (inputs(113));
    layer0_outputs(1419) <= not((inputs(139)) xor (inputs(189)));
    layer0_outputs(1420) <= not((inputs(59)) or (inputs(93)));
    layer0_outputs(1421) <= (inputs(49)) xor (inputs(227));
    layer0_outputs(1422) <= not(inputs(213));
    layer0_outputs(1423) <= inputs(212);
    layer0_outputs(1424) <= not(inputs(77));
    layer0_outputs(1425) <= not(inputs(172)) or (inputs(240));
    layer0_outputs(1426) <= (inputs(168)) and not (inputs(192));
    layer0_outputs(1427) <= inputs(55);
    layer0_outputs(1428) <= not(inputs(40)) or (inputs(94));
    layer0_outputs(1429) <= not((inputs(145)) and (inputs(72)));
    layer0_outputs(1430) <= not((inputs(82)) xor (inputs(217)));
    layer0_outputs(1431) <= not((inputs(7)) or (inputs(239)));
    layer0_outputs(1432) <= not((inputs(106)) or (inputs(54)));
    layer0_outputs(1433) <= inputs(232);
    layer0_outputs(1434) <= (inputs(146)) and not (inputs(27));
    layer0_outputs(1435) <= (inputs(123)) and not (inputs(104));
    layer0_outputs(1436) <= (inputs(3)) or (inputs(243));
    layer0_outputs(1437) <= not((inputs(67)) or (inputs(1)));
    layer0_outputs(1438) <= inputs(236);
    layer0_outputs(1439) <= not(inputs(73));
    layer0_outputs(1440) <= not((inputs(13)) and (inputs(249)));
    layer0_outputs(1441) <= not((inputs(169)) and (inputs(171)));
    layer0_outputs(1442) <= inputs(151);
    layer0_outputs(1443) <= '1';
    layer0_outputs(1444) <= not(inputs(123));
    layer0_outputs(1445) <= not(inputs(213)) or (inputs(109));
    layer0_outputs(1446) <= not((inputs(213)) or (inputs(128)));
    layer0_outputs(1447) <= inputs(180);
    layer0_outputs(1448) <= (inputs(216)) xor (inputs(247));
    layer0_outputs(1449) <= inputs(226);
    layer0_outputs(1450) <= (inputs(58)) or (inputs(3));
    layer0_outputs(1451) <= not(inputs(207)) or (inputs(230));
    layer0_outputs(1452) <= (inputs(22)) and not (inputs(251));
    layer0_outputs(1453) <= not((inputs(138)) and (inputs(106)));
    layer0_outputs(1454) <= inputs(83);
    layer0_outputs(1455) <= (inputs(170)) and not (inputs(41));
    layer0_outputs(1456) <= not((inputs(110)) xor (inputs(149)));
    layer0_outputs(1457) <= '1';
    layer0_outputs(1458) <= (inputs(161)) and not (inputs(28));
    layer0_outputs(1459) <= (inputs(59)) and (inputs(103));
    layer0_outputs(1460) <= inputs(241);
    layer0_outputs(1461) <= inputs(131);
    layer0_outputs(1462) <= not(inputs(84));
    layer0_outputs(1463) <= not(inputs(163));
    layer0_outputs(1464) <= not((inputs(25)) and (inputs(2)));
    layer0_outputs(1465) <= (inputs(238)) or (inputs(136));
    layer0_outputs(1466) <= (inputs(37)) and not (inputs(208));
    layer0_outputs(1467) <= (inputs(169)) xor (inputs(183));
    layer0_outputs(1468) <= (inputs(150)) and not (inputs(57));
    layer0_outputs(1469) <= (inputs(98)) or (inputs(162));
    layer0_outputs(1470) <= (inputs(135)) and not (inputs(170));
    layer0_outputs(1471) <= not(inputs(152));
    layer0_outputs(1472) <= inputs(2);
    layer0_outputs(1473) <= (inputs(166)) and not (inputs(143));
    layer0_outputs(1474) <= not(inputs(194));
    layer0_outputs(1475) <= not(inputs(7));
    layer0_outputs(1476) <= (inputs(148)) xor (inputs(105));
    layer0_outputs(1477) <= not(inputs(142)) or (inputs(224));
    layer0_outputs(1478) <= not((inputs(144)) or (inputs(143)));
    layer0_outputs(1479) <= '1';
    layer0_outputs(1480) <= not(inputs(50));
    layer0_outputs(1481) <= not((inputs(26)) or (inputs(248)));
    layer0_outputs(1482) <= not((inputs(241)) xor (inputs(247)));
    layer0_outputs(1483) <= not(inputs(25)) or (inputs(144));
    layer0_outputs(1484) <= not((inputs(39)) or (inputs(143)));
    layer0_outputs(1485) <= inputs(97);
    layer0_outputs(1486) <= (inputs(233)) xor (inputs(157));
    layer0_outputs(1487) <= not(inputs(19));
    layer0_outputs(1488) <= not((inputs(7)) or (inputs(203)));
    layer0_outputs(1489) <= not(inputs(179)) or (inputs(63));
    layer0_outputs(1490) <= not(inputs(184)) or (inputs(253));
    layer0_outputs(1491) <= inputs(75);
    layer0_outputs(1492) <= inputs(149);
    layer0_outputs(1493) <= (inputs(66)) and not (inputs(92));
    layer0_outputs(1494) <= (inputs(23)) and (inputs(26));
    layer0_outputs(1495) <= (inputs(127)) xor (inputs(136));
    layer0_outputs(1496) <= (inputs(136)) or (inputs(99));
    layer0_outputs(1497) <= (inputs(26)) and not (inputs(211));
    layer0_outputs(1498) <= not((inputs(91)) or (inputs(64)));
    layer0_outputs(1499) <= (inputs(189)) and not (inputs(248));
    layer0_outputs(1500) <= not((inputs(39)) or (inputs(24)));
    layer0_outputs(1501) <= inputs(250);
    layer0_outputs(1502) <= (inputs(12)) or (inputs(97));
    layer0_outputs(1503) <= not(inputs(139));
    layer0_outputs(1504) <= (inputs(8)) or (inputs(226));
    layer0_outputs(1505) <= not((inputs(230)) or (inputs(173)));
    layer0_outputs(1506) <= not(inputs(118));
    layer0_outputs(1507) <= not(inputs(46));
    layer0_outputs(1508) <= (inputs(103)) xor (inputs(207));
    layer0_outputs(1509) <= not(inputs(147)) or (inputs(33));
    layer0_outputs(1510) <= not(inputs(132));
    layer0_outputs(1511) <= not((inputs(64)) or (inputs(24)));
    layer0_outputs(1512) <= inputs(225);
    layer0_outputs(1513) <= (inputs(225)) and (inputs(222));
    layer0_outputs(1514) <= not((inputs(7)) xor (inputs(124)));
    layer0_outputs(1515) <= (inputs(230)) or (inputs(214));
    layer0_outputs(1516) <= (inputs(1)) or (inputs(127));
    layer0_outputs(1517) <= not(inputs(18)) or (inputs(151));
    layer0_outputs(1518) <= '0';
    layer0_outputs(1519) <= '0';
    layer0_outputs(1520) <= inputs(203);
    layer0_outputs(1521) <= not((inputs(183)) xor (inputs(35)));
    layer0_outputs(1522) <= not(inputs(93));
    layer0_outputs(1523) <= not((inputs(122)) or (inputs(47)));
    layer0_outputs(1524) <= not((inputs(46)) or (inputs(151)));
    layer0_outputs(1525) <= (inputs(129)) xor (inputs(101));
    layer0_outputs(1526) <= '1';
    layer0_outputs(1527) <= not(inputs(81)) or (inputs(110));
    layer0_outputs(1528) <= not((inputs(183)) xor (inputs(64)));
    layer0_outputs(1529) <= inputs(247);
    layer0_outputs(1530) <= not((inputs(84)) or (inputs(38)));
    layer0_outputs(1531) <= not(inputs(63)) or (inputs(215));
    layer0_outputs(1532) <= '1';
    layer0_outputs(1533) <= (inputs(179)) and (inputs(141));
    layer0_outputs(1534) <= (inputs(159)) xor (inputs(149));
    layer0_outputs(1535) <= '1';
    layer0_outputs(1536) <= (inputs(17)) xor (inputs(213));
    layer0_outputs(1537) <= not((inputs(216)) and (inputs(4)));
    layer0_outputs(1538) <= (inputs(197)) and not (inputs(251));
    layer0_outputs(1539) <= inputs(52);
    layer0_outputs(1540) <= (inputs(180)) and not (inputs(74));
    layer0_outputs(1541) <= inputs(17);
    layer0_outputs(1542) <= '1';
    layer0_outputs(1543) <= not((inputs(185)) xor (inputs(176)));
    layer0_outputs(1544) <= not((inputs(228)) and (inputs(14)));
    layer0_outputs(1545) <= inputs(231);
    layer0_outputs(1546) <= (inputs(243)) xor (inputs(232));
    layer0_outputs(1547) <= not((inputs(28)) and (inputs(234)));
    layer0_outputs(1548) <= (inputs(96)) or (inputs(128));
    layer0_outputs(1549) <= not(inputs(34));
    layer0_outputs(1550) <= not(inputs(203));
    layer0_outputs(1551) <= '0';
    layer0_outputs(1552) <= inputs(93);
    layer0_outputs(1553) <= not((inputs(233)) or (inputs(220)));
    layer0_outputs(1554) <= not((inputs(230)) or (inputs(192)));
    layer0_outputs(1555) <= not((inputs(124)) and (inputs(192)));
    layer0_outputs(1556) <= not(inputs(19));
    layer0_outputs(1557) <= (inputs(227)) and not (inputs(24));
    layer0_outputs(1558) <= '1';
    layer0_outputs(1559) <= not((inputs(161)) or (inputs(148)));
    layer0_outputs(1560) <= (inputs(50)) and not (inputs(60));
    layer0_outputs(1561) <= '1';
    layer0_outputs(1562) <= inputs(196);
    layer0_outputs(1563) <= '1';
    layer0_outputs(1564) <= (inputs(130)) or (inputs(92));
    layer0_outputs(1565) <= inputs(17);
    layer0_outputs(1566) <= inputs(178);
    layer0_outputs(1567) <= not(inputs(3)) or (inputs(175));
    layer0_outputs(1568) <= inputs(72);
    layer0_outputs(1569) <= not(inputs(165));
    layer0_outputs(1570) <= not(inputs(163)) or (inputs(190));
    layer0_outputs(1571) <= (inputs(48)) and not (inputs(114));
    layer0_outputs(1572) <= inputs(96);
    layer0_outputs(1573) <= not((inputs(71)) and (inputs(248)));
    layer0_outputs(1574) <= not(inputs(88));
    layer0_outputs(1575) <= (inputs(67)) and not (inputs(146));
    layer0_outputs(1576) <= not((inputs(117)) and (inputs(232)));
    layer0_outputs(1577) <= (inputs(246)) and not (inputs(16));
    layer0_outputs(1578) <= not((inputs(253)) or (inputs(2)));
    layer0_outputs(1579) <= inputs(145);
    layer0_outputs(1580) <= not((inputs(146)) or (inputs(144)));
    layer0_outputs(1581) <= not(inputs(217));
    layer0_outputs(1582) <= not(inputs(53)) or (inputs(123));
    layer0_outputs(1583) <= (inputs(138)) and not (inputs(224));
    layer0_outputs(1584) <= (inputs(206)) and (inputs(184));
    layer0_outputs(1585) <= '1';
    layer0_outputs(1586) <= not((inputs(102)) and (inputs(251)));
    layer0_outputs(1587) <= inputs(151);
    layer0_outputs(1588) <= (inputs(170)) and not (inputs(147));
    layer0_outputs(1589) <= inputs(115);
    layer0_outputs(1590) <= inputs(150);
    layer0_outputs(1591) <= not((inputs(140)) or (inputs(111)));
    layer0_outputs(1592) <= not((inputs(108)) xor (inputs(73)));
    layer0_outputs(1593) <= (inputs(62)) or (inputs(142));
    layer0_outputs(1594) <= inputs(194);
    layer0_outputs(1595) <= not((inputs(33)) or (inputs(21)));
    layer0_outputs(1596) <= not(inputs(37));
    layer0_outputs(1597) <= not((inputs(108)) xor (inputs(1)));
    layer0_outputs(1598) <= not(inputs(157));
    layer0_outputs(1599) <= not(inputs(86)) or (inputs(130));
    layer0_outputs(1600) <= not(inputs(160));
    layer0_outputs(1601) <= '1';
    layer0_outputs(1602) <= not(inputs(199)) or (inputs(217));
    layer0_outputs(1603) <= not(inputs(69));
    layer0_outputs(1604) <= not(inputs(121));
    layer0_outputs(1605) <= (inputs(62)) or (inputs(35));
    layer0_outputs(1606) <= not(inputs(72)) or (inputs(59));
    layer0_outputs(1607) <= not((inputs(139)) and (inputs(114)));
    layer0_outputs(1608) <= (inputs(26)) xor (inputs(160));
    layer0_outputs(1609) <= not((inputs(184)) or (inputs(87)));
    layer0_outputs(1610) <= not(inputs(163));
    layer0_outputs(1611) <= not(inputs(18)) or (inputs(163));
    layer0_outputs(1612) <= (inputs(215)) or (inputs(229));
    layer0_outputs(1613) <= not(inputs(74)) or (inputs(244));
    layer0_outputs(1614) <= not((inputs(27)) xor (inputs(62)));
    layer0_outputs(1615) <= not(inputs(241));
    layer0_outputs(1616) <= not((inputs(248)) xor (inputs(14)));
    layer0_outputs(1617) <= not((inputs(174)) or (inputs(249)));
    layer0_outputs(1618) <= not(inputs(154)) or (inputs(62));
    layer0_outputs(1619) <= inputs(78);
    layer0_outputs(1620) <= not(inputs(116));
    layer0_outputs(1621) <= (inputs(13)) xor (inputs(6));
    layer0_outputs(1622) <= inputs(48);
    layer0_outputs(1623) <= not(inputs(21));
    layer0_outputs(1624) <= '0';
    layer0_outputs(1625) <= inputs(90);
    layer0_outputs(1626) <= (inputs(62)) and (inputs(196));
    layer0_outputs(1627) <= (inputs(166)) and not (inputs(191));
    layer0_outputs(1628) <= not(inputs(164));
    layer0_outputs(1629) <= (inputs(59)) and not (inputs(21));
    layer0_outputs(1630) <= not((inputs(44)) or (inputs(17)));
    layer0_outputs(1631) <= not(inputs(231));
    layer0_outputs(1632) <= not(inputs(108));
    layer0_outputs(1633) <= not((inputs(201)) and (inputs(173)));
    layer0_outputs(1634) <= '0';
    layer0_outputs(1635) <= not(inputs(98)) or (inputs(243));
    layer0_outputs(1636) <= not(inputs(105));
    layer0_outputs(1637) <= inputs(3);
    layer0_outputs(1638) <= not((inputs(7)) or (inputs(3)));
    layer0_outputs(1639) <= not((inputs(10)) xor (inputs(96)));
    layer0_outputs(1640) <= (inputs(9)) or (inputs(61));
    layer0_outputs(1641) <= '0';
    layer0_outputs(1642) <= not(inputs(26)) or (inputs(175));
    layer0_outputs(1643) <= (inputs(139)) and not (inputs(250));
    layer0_outputs(1644) <= not((inputs(67)) or (inputs(166)));
    layer0_outputs(1645) <= inputs(167);
    layer0_outputs(1646) <= inputs(23);
    layer0_outputs(1647) <= '0';
    layer0_outputs(1648) <= (inputs(179)) and not (inputs(102));
    layer0_outputs(1649) <= (inputs(83)) xor (inputs(111));
    layer0_outputs(1650) <= not((inputs(77)) xor (inputs(41)));
    layer0_outputs(1651) <= inputs(128);
    layer0_outputs(1652) <= not((inputs(222)) or (inputs(206)));
    layer0_outputs(1653) <= not((inputs(218)) or (inputs(125)));
    layer0_outputs(1654) <= (inputs(70)) and (inputs(101));
    layer0_outputs(1655) <= not((inputs(34)) xor (inputs(79)));
    layer0_outputs(1656) <= (inputs(223)) or (inputs(22));
    layer0_outputs(1657) <= not((inputs(225)) or (inputs(81)));
    layer0_outputs(1658) <= '1';
    layer0_outputs(1659) <= (inputs(176)) and not (inputs(207));
    layer0_outputs(1660) <= not((inputs(96)) or (inputs(245)));
    layer0_outputs(1661) <= not(inputs(195)) or (inputs(239));
    layer0_outputs(1662) <= not(inputs(75)) or (inputs(147));
    layer0_outputs(1663) <= not(inputs(150));
    layer0_outputs(1664) <= (inputs(84)) and not (inputs(87));
    layer0_outputs(1665) <= inputs(103);
    layer0_outputs(1666) <= not(inputs(41));
    layer0_outputs(1667) <= not((inputs(194)) xor (inputs(242)));
    layer0_outputs(1668) <= (inputs(121)) or (inputs(110));
    layer0_outputs(1669) <= (inputs(80)) or (inputs(94));
    layer0_outputs(1670) <= (inputs(120)) xor (inputs(134));
    layer0_outputs(1671) <= not((inputs(92)) xor (inputs(106)));
    layer0_outputs(1672) <= not(inputs(101)) or (inputs(94));
    layer0_outputs(1673) <= not(inputs(65)) or (inputs(145));
    layer0_outputs(1674) <= (inputs(31)) and not (inputs(169));
    layer0_outputs(1675) <= not((inputs(30)) xor (inputs(4)));
    layer0_outputs(1676) <= (inputs(13)) xor (inputs(206));
    layer0_outputs(1677) <= not(inputs(18));
    layer0_outputs(1678) <= '1';
    layer0_outputs(1679) <= (inputs(71)) and not (inputs(32));
    layer0_outputs(1680) <= not(inputs(0)) or (inputs(50));
    layer0_outputs(1681) <= not(inputs(91)) or (inputs(227));
    layer0_outputs(1682) <= (inputs(131)) and not (inputs(117));
    layer0_outputs(1683) <= not(inputs(249)) or (inputs(227));
    layer0_outputs(1684) <= not(inputs(7)) or (inputs(177));
    layer0_outputs(1685) <= inputs(148);
    layer0_outputs(1686) <= not(inputs(78)) or (inputs(220));
    layer0_outputs(1687) <= (inputs(186)) or (inputs(142));
    layer0_outputs(1688) <= not(inputs(84));
    layer0_outputs(1689) <= not(inputs(119));
    layer0_outputs(1690) <= '0';
    layer0_outputs(1691) <= not((inputs(218)) or (inputs(157)));
    layer0_outputs(1692) <= not(inputs(167)) or (inputs(208));
    layer0_outputs(1693) <= (inputs(149)) xor (inputs(14));
    layer0_outputs(1694) <= not(inputs(68)) or (inputs(220));
    layer0_outputs(1695) <= inputs(91);
    layer0_outputs(1696) <= not(inputs(103)) or (inputs(18));
    layer0_outputs(1697) <= inputs(135);
    layer0_outputs(1698) <= (inputs(166)) and not (inputs(248));
    layer0_outputs(1699) <= not(inputs(20)) or (inputs(142));
    layer0_outputs(1700) <= not((inputs(173)) or (inputs(72)));
    layer0_outputs(1701) <= not((inputs(166)) xor (inputs(123)));
    layer0_outputs(1702) <= not((inputs(116)) or (inputs(80)));
    layer0_outputs(1703) <= (inputs(199)) and not (inputs(107));
    layer0_outputs(1704) <= not((inputs(105)) xor (inputs(187)));
    layer0_outputs(1705) <= not(inputs(166)) or (inputs(146));
    layer0_outputs(1706) <= (inputs(255)) xor (inputs(89));
    layer0_outputs(1707) <= (inputs(17)) and not (inputs(82));
    layer0_outputs(1708) <= inputs(168);
    layer0_outputs(1709) <= '1';
    layer0_outputs(1710) <= '1';
    layer0_outputs(1711) <= not(inputs(100));
    layer0_outputs(1712) <= (inputs(134)) or (inputs(41));
    layer0_outputs(1713) <= (inputs(74)) or (inputs(88));
    layer0_outputs(1714) <= not(inputs(172));
    layer0_outputs(1715) <= not(inputs(196));
    layer0_outputs(1716) <= not((inputs(178)) xor (inputs(252)));
    layer0_outputs(1717) <= (inputs(116)) and not (inputs(207));
    layer0_outputs(1718) <= (inputs(78)) or (inputs(174));
    layer0_outputs(1719) <= not(inputs(188)) or (inputs(15));
    layer0_outputs(1720) <= not((inputs(236)) or (inputs(121)));
    layer0_outputs(1721) <= not((inputs(244)) and (inputs(104)));
    layer0_outputs(1722) <= (inputs(138)) xor (inputs(103));
    layer0_outputs(1723) <= not(inputs(130));
    layer0_outputs(1724) <= (inputs(160)) and (inputs(160));
    layer0_outputs(1725) <= not(inputs(19)) or (inputs(4));
    layer0_outputs(1726) <= (inputs(229)) or (inputs(227));
    layer0_outputs(1727) <= (inputs(191)) and not (inputs(107));
    layer0_outputs(1728) <= not(inputs(141)) or (inputs(13));
    layer0_outputs(1729) <= not(inputs(198));
    layer0_outputs(1730) <= (inputs(147)) or (inputs(148));
    layer0_outputs(1731) <= (inputs(79)) xor (inputs(28));
    layer0_outputs(1732) <= (inputs(60)) or (inputs(19));
    layer0_outputs(1733) <= not((inputs(211)) or (inputs(212)));
    layer0_outputs(1734) <= not(inputs(136)) or (inputs(187));
    layer0_outputs(1735) <= not(inputs(30));
    layer0_outputs(1736) <= inputs(118);
    layer0_outputs(1737) <= (inputs(72)) xor (inputs(45));
    layer0_outputs(1738) <= (inputs(21)) or (inputs(94));
    layer0_outputs(1739) <= (inputs(28)) xor (inputs(42));
    layer0_outputs(1740) <= not(inputs(143));
    layer0_outputs(1741) <= not((inputs(72)) xor (inputs(171)));
    layer0_outputs(1742) <= inputs(67);
    layer0_outputs(1743) <= not((inputs(128)) xor (inputs(205)));
    layer0_outputs(1744) <= not(inputs(172)) or (inputs(184));
    layer0_outputs(1745) <= inputs(97);
    layer0_outputs(1746) <= not(inputs(203));
    layer0_outputs(1747) <= not(inputs(62)) or (inputs(249));
    layer0_outputs(1748) <= (inputs(212)) and not (inputs(117));
    layer0_outputs(1749) <= (inputs(83)) and not (inputs(209));
    layer0_outputs(1750) <= not((inputs(109)) and (inputs(237)));
    layer0_outputs(1751) <= not((inputs(250)) or (inputs(233)));
    layer0_outputs(1752) <= not(inputs(191));
    layer0_outputs(1753) <= not((inputs(117)) or (inputs(170)));
    layer0_outputs(1754) <= inputs(30);
    layer0_outputs(1755) <= not(inputs(90)) or (inputs(190));
    layer0_outputs(1756) <= not(inputs(254)) or (inputs(191));
    layer0_outputs(1757) <= (inputs(25)) and not (inputs(203));
    layer0_outputs(1758) <= not(inputs(194));
    layer0_outputs(1759) <= not(inputs(212)) or (inputs(134));
    layer0_outputs(1760) <= (inputs(197)) and not (inputs(91));
    layer0_outputs(1761) <= not(inputs(158));
    layer0_outputs(1762) <= inputs(145);
    layer0_outputs(1763) <= not((inputs(77)) or (inputs(150)));
    layer0_outputs(1764) <= '0';
    layer0_outputs(1765) <= not((inputs(119)) or (inputs(20)));
    layer0_outputs(1766) <= (inputs(208)) or (inputs(114));
    layer0_outputs(1767) <= not((inputs(138)) or (inputs(202)));
    layer0_outputs(1768) <= (inputs(186)) and (inputs(122));
    layer0_outputs(1769) <= '1';
    layer0_outputs(1770) <= not(inputs(88));
    layer0_outputs(1771) <= not(inputs(234));
    layer0_outputs(1772) <= inputs(79);
    layer0_outputs(1773) <= inputs(152);
    layer0_outputs(1774) <= not(inputs(34));
    layer0_outputs(1775) <= not(inputs(147)) or (inputs(211));
    layer0_outputs(1776) <= (inputs(208)) or (inputs(116));
    layer0_outputs(1777) <= not(inputs(151));
    layer0_outputs(1778) <= not((inputs(69)) or (inputs(165)));
    layer0_outputs(1779) <= not((inputs(46)) and (inputs(118)));
    layer0_outputs(1780) <= inputs(79);
    layer0_outputs(1781) <= not((inputs(233)) or (inputs(131)));
    layer0_outputs(1782) <= inputs(57);
    layer0_outputs(1783) <= not((inputs(61)) xor (inputs(230)));
    layer0_outputs(1784) <= not((inputs(205)) or (inputs(88)));
    layer0_outputs(1785) <= not(inputs(77));
    layer0_outputs(1786) <= not(inputs(105));
    layer0_outputs(1787) <= inputs(203);
    layer0_outputs(1788) <= (inputs(38)) and not (inputs(190));
    layer0_outputs(1789) <= '1';
    layer0_outputs(1790) <= not((inputs(66)) and (inputs(161)));
    layer0_outputs(1791) <= (inputs(170)) or (inputs(43));
    layer0_outputs(1792) <= not(inputs(34)) or (inputs(39));
    layer0_outputs(1793) <= inputs(173);
    layer0_outputs(1794) <= (inputs(17)) or (inputs(44));
    layer0_outputs(1795) <= '0';
    layer0_outputs(1796) <= not(inputs(168)) or (inputs(60));
    layer0_outputs(1797) <= not(inputs(16)) or (inputs(238));
    layer0_outputs(1798) <= not((inputs(152)) or (inputs(16)));
    layer0_outputs(1799) <= not((inputs(93)) or (inputs(79)));
    layer0_outputs(1800) <= not(inputs(173));
    layer0_outputs(1801) <= not((inputs(43)) xor (inputs(92)));
    layer0_outputs(1802) <= not(inputs(90)) or (inputs(56));
    layer0_outputs(1803) <= not(inputs(200)) or (inputs(89));
    layer0_outputs(1804) <= (inputs(52)) xor (inputs(4));
    layer0_outputs(1805) <= (inputs(114)) and not (inputs(241));
    layer0_outputs(1806) <= (inputs(160)) and not (inputs(175));
    layer0_outputs(1807) <= not((inputs(236)) or (inputs(197)));
    layer0_outputs(1808) <= not(inputs(10));
    layer0_outputs(1809) <= not((inputs(62)) or (inputs(63)));
    layer0_outputs(1810) <= (inputs(145)) xor (inputs(164));
    layer0_outputs(1811) <= (inputs(53)) and not (inputs(172));
    layer0_outputs(1812) <= not(inputs(151));
    layer0_outputs(1813) <= not(inputs(247));
    layer0_outputs(1814) <= inputs(160);
    layer0_outputs(1815) <= not((inputs(232)) and (inputs(213)));
    layer0_outputs(1816) <= (inputs(109)) or (inputs(165));
    layer0_outputs(1817) <= (inputs(46)) xor (inputs(74));
    layer0_outputs(1818) <= '1';
    layer0_outputs(1819) <= inputs(176);
    layer0_outputs(1820) <= not((inputs(181)) xor (inputs(227)));
    layer0_outputs(1821) <= inputs(174);
    layer0_outputs(1822) <= not(inputs(198)) or (inputs(174));
    layer0_outputs(1823) <= inputs(58);
    layer0_outputs(1824) <= (inputs(162)) and not (inputs(113));
    layer0_outputs(1825) <= inputs(0);
    layer0_outputs(1826) <= inputs(45);
    layer0_outputs(1827) <= (inputs(63)) or (inputs(250));
    layer0_outputs(1828) <= not(inputs(5));
    layer0_outputs(1829) <= (inputs(6)) xor (inputs(53));
    layer0_outputs(1830) <= not(inputs(100)) or (inputs(159));
    layer0_outputs(1831) <= not(inputs(137)) or (inputs(176));
    layer0_outputs(1832) <= (inputs(88)) xor (inputs(112));
    layer0_outputs(1833) <= (inputs(209)) or (inputs(244));
    layer0_outputs(1834) <= not(inputs(180)) or (inputs(252));
    layer0_outputs(1835) <= not((inputs(2)) or (inputs(0)));
    layer0_outputs(1836) <= inputs(179);
    layer0_outputs(1837) <= not(inputs(86));
    layer0_outputs(1838) <= not(inputs(210)) or (inputs(71));
    layer0_outputs(1839) <= inputs(190);
    layer0_outputs(1840) <= not((inputs(12)) or (inputs(65)));
    layer0_outputs(1841) <= (inputs(79)) and (inputs(238));
    layer0_outputs(1842) <= inputs(22);
    layer0_outputs(1843) <= inputs(202);
    layer0_outputs(1844) <= (inputs(243)) and not (inputs(97));
    layer0_outputs(1845) <= (inputs(174)) xor (inputs(165));
    layer0_outputs(1846) <= not((inputs(112)) or (inputs(212)));
    layer0_outputs(1847) <= not(inputs(134)) or (inputs(33));
    layer0_outputs(1848) <= not((inputs(211)) xor (inputs(212)));
    layer0_outputs(1849) <= (inputs(233)) and not (inputs(156));
    layer0_outputs(1850) <= not(inputs(100));
    layer0_outputs(1851) <= not(inputs(48));
    layer0_outputs(1852) <= (inputs(163)) or (inputs(111));
    layer0_outputs(1853) <= not(inputs(136)) or (inputs(53));
    layer0_outputs(1854) <= not(inputs(245));
    layer0_outputs(1855) <= not(inputs(181));
    layer0_outputs(1856) <= inputs(86);
    layer0_outputs(1857) <= not((inputs(130)) or (inputs(227)));
    layer0_outputs(1858) <= (inputs(44)) or (inputs(38));
    layer0_outputs(1859) <= not(inputs(187));
    layer0_outputs(1860) <= not(inputs(22)) or (inputs(146));
    layer0_outputs(1861) <= not(inputs(165));
    layer0_outputs(1862) <= not((inputs(228)) or (inputs(30)));
    layer0_outputs(1863) <= not(inputs(231));
    layer0_outputs(1864) <= '0';
    layer0_outputs(1865) <= not(inputs(212));
    layer0_outputs(1866) <= (inputs(174)) or (inputs(219));
    layer0_outputs(1867) <= (inputs(243)) and not (inputs(70));
    layer0_outputs(1868) <= inputs(79);
    layer0_outputs(1869) <= not(inputs(27)) or (inputs(188));
    layer0_outputs(1870) <= not(inputs(213));
    layer0_outputs(1871) <= (inputs(17)) and not (inputs(14));
    layer0_outputs(1872) <= not(inputs(109));
    layer0_outputs(1873) <= not(inputs(58)) or (inputs(152));
    layer0_outputs(1874) <= inputs(146);
    layer0_outputs(1875) <= not((inputs(218)) or (inputs(191)));
    layer0_outputs(1876) <= (inputs(27)) and (inputs(228));
    layer0_outputs(1877) <= inputs(4);
    layer0_outputs(1878) <= not((inputs(82)) xor (inputs(85)));
    layer0_outputs(1879) <= inputs(21);
    layer0_outputs(1880) <= not(inputs(178)) or (inputs(113));
    layer0_outputs(1881) <= (inputs(109)) or (inputs(36));
    layer0_outputs(1882) <= not((inputs(169)) or (inputs(167)));
    layer0_outputs(1883) <= not((inputs(71)) xor (inputs(192)));
    layer0_outputs(1884) <= inputs(4);
    layer0_outputs(1885) <= not(inputs(51)) or (inputs(213));
    layer0_outputs(1886) <= (inputs(68)) or (inputs(142));
    layer0_outputs(1887) <= not((inputs(194)) or (inputs(252)));
    layer0_outputs(1888) <= not(inputs(218)) or (inputs(177));
    layer0_outputs(1889) <= inputs(85);
    layer0_outputs(1890) <= not((inputs(201)) and (inputs(238)));
    layer0_outputs(1891) <= not(inputs(118));
    layer0_outputs(1892) <= (inputs(9)) and (inputs(28));
    layer0_outputs(1893) <= inputs(247);
    layer0_outputs(1894) <= not(inputs(216));
    layer0_outputs(1895) <= inputs(46);
    layer0_outputs(1896) <= (inputs(41)) and not (inputs(255));
    layer0_outputs(1897) <= not(inputs(202)) or (inputs(242));
    layer0_outputs(1898) <= (inputs(172)) xor (inputs(60));
    layer0_outputs(1899) <= not(inputs(193));
    layer0_outputs(1900) <= (inputs(100)) and not (inputs(66));
    layer0_outputs(1901) <= not(inputs(165));
    layer0_outputs(1902) <= not(inputs(93));
    layer0_outputs(1903) <= inputs(233);
    layer0_outputs(1904) <= not(inputs(191));
    layer0_outputs(1905) <= inputs(228);
    layer0_outputs(1906) <= not(inputs(140)) or (inputs(48));
    layer0_outputs(1907) <= not(inputs(114));
    layer0_outputs(1908) <= not(inputs(81)) or (inputs(184));
    layer0_outputs(1909) <= not((inputs(253)) xor (inputs(139)));
    layer0_outputs(1910) <= not((inputs(76)) or (inputs(238)));
    layer0_outputs(1911) <= (inputs(219)) xor (inputs(156));
    layer0_outputs(1912) <= not(inputs(165));
    layer0_outputs(1913) <= (inputs(246)) and not (inputs(36));
    layer0_outputs(1914) <= inputs(239);
    layer0_outputs(1915) <= inputs(88);
    layer0_outputs(1916) <= (inputs(187)) or (inputs(26));
    layer0_outputs(1917) <= inputs(162);
    layer0_outputs(1918) <= not((inputs(116)) or (inputs(175)));
    layer0_outputs(1919) <= inputs(158);
    layer0_outputs(1920) <= not(inputs(210));
    layer0_outputs(1921) <= not(inputs(164));
    layer0_outputs(1922) <= inputs(88);
    layer0_outputs(1923) <= not(inputs(246));
    layer0_outputs(1924) <= '1';
    layer0_outputs(1925) <= inputs(59);
    layer0_outputs(1926) <= not(inputs(165)) or (inputs(0));
    layer0_outputs(1927) <= not(inputs(44)) or (inputs(252));
    layer0_outputs(1928) <= not(inputs(38)) or (inputs(195));
    layer0_outputs(1929) <= not((inputs(200)) or (inputs(40)));
    layer0_outputs(1930) <= inputs(231);
    layer0_outputs(1931) <= not((inputs(226)) and (inputs(6)));
    layer0_outputs(1932) <= not(inputs(195));
    layer0_outputs(1933) <= (inputs(82)) or (inputs(50));
    layer0_outputs(1934) <= inputs(124);
    layer0_outputs(1935) <= (inputs(14)) and (inputs(15));
    layer0_outputs(1936) <= (inputs(120)) or (inputs(6));
    layer0_outputs(1937) <= not((inputs(159)) or (inputs(102)));
    layer0_outputs(1938) <= (inputs(27)) and not (inputs(143));
    layer0_outputs(1939) <= not((inputs(94)) xor (inputs(28)));
    layer0_outputs(1940) <= (inputs(83)) or (inputs(171));
    layer0_outputs(1941) <= not((inputs(91)) xor (inputs(18)));
    layer0_outputs(1942) <= not(inputs(144));
    layer0_outputs(1943) <= (inputs(79)) xor (inputs(91));
    layer0_outputs(1944) <= inputs(149);
    layer0_outputs(1945) <= not((inputs(53)) or (inputs(27)));
    layer0_outputs(1946) <= '0';
    layer0_outputs(1947) <= (inputs(190)) xor (inputs(113));
    layer0_outputs(1948) <= inputs(91);
    layer0_outputs(1949) <= not(inputs(134));
    layer0_outputs(1950) <= inputs(156);
    layer0_outputs(1951) <= not(inputs(17));
    layer0_outputs(1952) <= (inputs(80)) and (inputs(244));
    layer0_outputs(1953) <= (inputs(110)) and not (inputs(153));
    layer0_outputs(1954) <= inputs(69);
    layer0_outputs(1955) <= (inputs(192)) and not (inputs(253));
    layer0_outputs(1956) <= (inputs(104)) and not (inputs(236));
    layer0_outputs(1957) <= not(inputs(255));
    layer0_outputs(1958) <= inputs(96);
    layer0_outputs(1959) <= (inputs(243)) or (inputs(6));
    layer0_outputs(1960) <= not(inputs(200)) or (inputs(97));
    layer0_outputs(1961) <= (inputs(113)) and not (inputs(155));
    layer0_outputs(1962) <= inputs(254);
    layer0_outputs(1963) <= (inputs(125)) and (inputs(200));
    layer0_outputs(1964) <= (inputs(69)) xor (inputs(81));
    layer0_outputs(1965) <= inputs(81);
    layer0_outputs(1966) <= inputs(191);
    layer0_outputs(1967) <= not((inputs(99)) and (inputs(41)));
    layer0_outputs(1968) <= inputs(133);
    layer0_outputs(1969) <= not(inputs(18)) or (inputs(127));
    layer0_outputs(1970) <= not(inputs(99));
    layer0_outputs(1971) <= not(inputs(136)) or (inputs(115));
    layer0_outputs(1972) <= not(inputs(193));
    layer0_outputs(1973) <= inputs(114);
    layer0_outputs(1974) <= (inputs(231)) and not (inputs(207));
    layer0_outputs(1975) <= (inputs(65)) or (inputs(204));
    layer0_outputs(1976) <= '1';
    layer0_outputs(1977) <= not((inputs(36)) xor (inputs(166)));
    layer0_outputs(1978) <= not((inputs(72)) and (inputs(21)));
    layer0_outputs(1979) <= (inputs(191)) or (inputs(161));
    layer0_outputs(1980) <= (inputs(44)) and not (inputs(230));
    layer0_outputs(1981) <= not(inputs(11));
    layer0_outputs(1982) <= not(inputs(77));
    layer0_outputs(1983) <= not((inputs(66)) and (inputs(47)));
    layer0_outputs(1984) <= inputs(148);
    layer0_outputs(1985) <= not(inputs(136));
    layer0_outputs(1986) <= (inputs(130)) and not (inputs(155));
    layer0_outputs(1987) <= inputs(164);
    layer0_outputs(1988) <= not(inputs(62));
    layer0_outputs(1989) <= not((inputs(129)) xor (inputs(175)));
    layer0_outputs(1990) <= inputs(104);
    layer0_outputs(1991) <= (inputs(101)) and (inputs(79));
    layer0_outputs(1992) <= not((inputs(218)) or (inputs(185)));
    layer0_outputs(1993) <= '0';
    layer0_outputs(1994) <= not(inputs(150));
    layer0_outputs(1995) <= not((inputs(126)) or (inputs(188)));
    layer0_outputs(1996) <= inputs(99);
    layer0_outputs(1997) <= (inputs(226)) or (inputs(41));
    layer0_outputs(1998) <= (inputs(72)) xor (inputs(24));
    layer0_outputs(1999) <= (inputs(150)) or (inputs(227));
    layer0_outputs(2000) <= not((inputs(22)) or (inputs(5)));
    layer0_outputs(2001) <= inputs(250);
    layer0_outputs(2002) <= (inputs(18)) and not (inputs(144));
    layer0_outputs(2003) <= not((inputs(116)) and (inputs(200)));
    layer0_outputs(2004) <= not(inputs(190)) or (inputs(46));
    layer0_outputs(2005) <= (inputs(213)) and not (inputs(37));
    layer0_outputs(2006) <= not((inputs(147)) or (inputs(84)));
    layer0_outputs(2007) <= not(inputs(122));
    layer0_outputs(2008) <= not(inputs(182));
    layer0_outputs(2009) <= (inputs(179)) and not (inputs(157));
    layer0_outputs(2010) <= not((inputs(62)) xor (inputs(236)));
    layer0_outputs(2011) <= not(inputs(162));
    layer0_outputs(2012) <= not(inputs(85)) or (inputs(186));
    layer0_outputs(2013) <= (inputs(198)) and not (inputs(38));
    layer0_outputs(2014) <= not(inputs(105));
    layer0_outputs(2015) <= not((inputs(253)) or (inputs(137)));
    layer0_outputs(2016) <= not((inputs(53)) or (inputs(81)));
    layer0_outputs(2017) <= inputs(107);
    layer0_outputs(2018) <= not(inputs(6)) or (inputs(230));
    layer0_outputs(2019) <= (inputs(236)) or (inputs(81));
    layer0_outputs(2020) <= (inputs(44)) or (inputs(141));
    layer0_outputs(2021) <= not(inputs(29));
    layer0_outputs(2022) <= '1';
    layer0_outputs(2023) <= inputs(77);
    layer0_outputs(2024) <= not(inputs(103));
    layer0_outputs(2025) <= not(inputs(18));
    layer0_outputs(2026) <= inputs(183);
    layer0_outputs(2027) <= inputs(192);
    layer0_outputs(2028) <= (inputs(164)) and not (inputs(55));
    layer0_outputs(2029) <= inputs(56);
    layer0_outputs(2030) <= (inputs(140)) or (inputs(113));
    layer0_outputs(2031) <= (inputs(13)) and (inputs(13));
    layer0_outputs(2032) <= not((inputs(38)) and (inputs(74)));
    layer0_outputs(2033) <= not((inputs(26)) or (inputs(39)));
    layer0_outputs(2034) <= not((inputs(159)) or (inputs(219)));
    layer0_outputs(2035) <= inputs(230);
    layer0_outputs(2036) <= not((inputs(146)) or (inputs(126)));
    layer0_outputs(2037) <= (inputs(20)) and not (inputs(156));
    layer0_outputs(2038) <= not(inputs(237));
    layer0_outputs(2039) <= not(inputs(82));
    layer0_outputs(2040) <= inputs(251);
    layer0_outputs(2041) <= (inputs(17)) or (inputs(238));
    layer0_outputs(2042) <= not(inputs(22));
    layer0_outputs(2043) <= inputs(119);
    layer0_outputs(2044) <= not(inputs(142)) or (inputs(127));
    layer0_outputs(2045) <= inputs(88);
    layer0_outputs(2046) <= (inputs(164)) and not (inputs(78));
    layer0_outputs(2047) <= not((inputs(134)) or (inputs(160)));
    layer0_outputs(2048) <= inputs(177);
    layer0_outputs(2049) <= '0';
    layer0_outputs(2050) <= not(inputs(95));
    layer0_outputs(2051) <= not((inputs(89)) or (inputs(191)));
    layer0_outputs(2052) <= not((inputs(37)) or (inputs(125)));
    layer0_outputs(2053) <= '1';
    layer0_outputs(2054) <= not((inputs(70)) xor (inputs(183)));
    layer0_outputs(2055) <= (inputs(72)) xor (inputs(11));
    layer0_outputs(2056) <= (inputs(245)) or (inputs(98));
    layer0_outputs(2057) <= not((inputs(93)) or (inputs(7)));
    layer0_outputs(2058) <= not(inputs(107));
    layer0_outputs(2059) <= not(inputs(205));
    layer0_outputs(2060) <= not(inputs(166));
    layer0_outputs(2061) <= not(inputs(203));
    layer0_outputs(2062) <= (inputs(66)) or (inputs(205));
    layer0_outputs(2063) <= (inputs(216)) and (inputs(197));
    layer0_outputs(2064) <= not((inputs(43)) or (inputs(56)));
    layer0_outputs(2065) <= inputs(45);
    layer0_outputs(2066) <= not(inputs(229)) or (inputs(151));
    layer0_outputs(2067) <= not((inputs(154)) and (inputs(202)));
    layer0_outputs(2068) <= (inputs(176)) xor (inputs(186));
    layer0_outputs(2069) <= (inputs(125)) or (inputs(31));
    layer0_outputs(2070) <= not((inputs(54)) and (inputs(100)));
    layer0_outputs(2071) <= not((inputs(42)) xor (inputs(72)));
    layer0_outputs(2072) <= inputs(76);
    layer0_outputs(2073) <= not((inputs(178)) xor (inputs(126)));
    layer0_outputs(2074) <= not((inputs(235)) or (inputs(204)));
    layer0_outputs(2075) <= (inputs(88)) and not (inputs(54));
    layer0_outputs(2076) <= not(inputs(18)) or (inputs(11));
    layer0_outputs(2077) <= not((inputs(217)) or (inputs(233)));
    layer0_outputs(2078) <= inputs(25);
    layer0_outputs(2079) <= not(inputs(87));
    layer0_outputs(2080) <= not((inputs(178)) and (inputs(254)));
    layer0_outputs(2081) <= (inputs(34)) or (inputs(166));
    layer0_outputs(2082) <= not(inputs(154));
    layer0_outputs(2083) <= (inputs(118)) and not (inputs(8));
    layer0_outputs(2084) <= not(inputs(88));
    layer0_outputs(2085) <= (inputs(201)) xor (inputs(185));
    layer0_outputs(2086) <= not(inputs(155)) or (inputs(68));
    layer0_outputs(2087) <= (inputs(69)) xor (inputs(35));
    layer0_outputs(2088) <= not((inputs(40)) xor (inputs(157)));
    layer0_outputs(2089) <= (inputs(170)) and not (inputs(103));
    layer0_outputs(2090) <= (inputs(234)) or (inputs(35));
    layer0_outputs(2091) <= not(inputs(31));
    layer0_outputs(2092) <= not((inputs(112)) xor (inputs(129)));
    layer0_outputs(2093) <= not((inputs(208)) xor (inputs(150)));
    layer0_outputs(2094) <= not(inputs(36)) or (inputs(221));
    layer0_outputs(2095) <= not(inputs(98));
    layer0_outputs(2096) <= not((inputs(20)) or (inputs(25)));
    layer0_outputs(2097) <= not(inputs(136));
    layer0_outputs(2098) <= (inputs(186)) or (inputs(115));
    layer0_outputs(2099) <= not(inputs(121)) or (inputs(143));
    layer0_outputs(2100) <= not(inputs(250)) or (inputs(240));
    layer0_outputs(2101) <= not(inputs(221)) or (inputs(141));
    layer0_outputs(2102) <= (inputs(59)) and not (inputs(9));
    layer0_outputs(2103) <= (inputs(63)) xor (inputs(121));
    layer0_outputs(2104) <= inputs(131);
    layer0_outputs(2105) <= (inputs(8)) and not (inputs(18));
    layer0_outputs(2106) <= inputs(163);
    layer0_outputs(2107) <= inputs(39);
    layer0_outputs(2108) <= '0';
    layer0_outputs(2109) <= inputs(220);
    layer0_outputs(2110) <= not((inputs(189)) or (inputs(134)));
    layer0_outputs(2111) <= (inputs(36)) and (inputs(225));
    layer0_outputs(2112) <= (inputs(158)) and not (inputs(235));
    layer0_outputs(2113) <= inputs(196);
    layer0_outputs(2114) <= not((inputs(42)) or (inputs(31)));
    layer0_outputs(2115) <= not(inputs(156)) or (inputs(220));
    layer0_outputs(2116) <= not(inputs(137));
    layer0_outputs(2117) <= not(inputs(177));
    layer0_outputs(2118) <= not(inputs(167)) or (inputs(3));
    layer0_outputs(2119) <= not((inputs(200)) and (inputs(212)));
    layer0_outputs(2120) <= inputs(111);
    layer0_outputs(2121) <= not((inputs(61)) xor (inputs(253)));
    layer0_outputs(2122) <= not(inputs(57));
    layer0_outputs(2123) <= inputs(219);
    layer0_outputs(2124) <= not(inputs(93)) or (inputs(240));
    layer0_outputs(2125) <= (inputs(95)) and not (inputs(223));
    layer0_outputs(2126) <= inputs(38);
    layer0_outputs(2127) <= not((inputs(177)) xor (inputs(204)));
    layer0_outputs(2128) <= (inputs(49)) xor (inputs(204));
    layer0_outputs(2129) <= not(inputs(27));
    layer0_outputs(2130) <= not((inputs(209)) or (inputs(190)));
    layer0_outputs(2131) <= not(inputs(204));
    layer0_outputs(2132) <= not(inputs(205)) or (inputs(240));
    layer0_outputs(2133) <= (inputs(68)) xor (inputs(22));
    layer0_outputs(2134) <= (inputs(251)) and (inputs(65));
    layer0_outputs(2135) <= not(inputs(228));
    layer0_outputs(2136) <= (inputs(97)) or (inputs(30));
    layer0_outputs(2137) <= (inputs(99)) and not (inputs(217));
    layer0_outputs(2138) <= (inputs(198)) and not (inputs(95));
    layer0_outputs(2139) <= inputs(116);
    layer0_outputs(2140) <= '0';
    layer0_outputs(2141) <= (inputs(57)) and not (inputs(255));
    layer0_outputs(2142) <= inputs(99);
    layer0_outputs(2143) <= inputs(108);
    layer0_outputs(2144) <= inputs(230);
    layer0_outputs(2145) <= not((inputs(124)) or (inputs(20)));
    layer0_outputs(2146) <= (inputs(110)) xor (inputs(22));
    layer0_outputs(2147) <= not((inputs(54)) xor (inputs(249)));
    layer0_outputs(2148) <= (inputs(121)) and not (inputs(114));
    layer0_outputs(2149) <= (inputs(121)) and not (inputs(10));
    layer0_outputs(2150) <= not((inputs(3)) and (inputs(155)));
    layer0_outputs(2151) <= (inputs(39)) or (inputs(174));
    layer0_outputs(2152) <= inputs(114);
    layer0_outputs(2153) <= (inputs(53)) and not (inputs(191));
    layer0_outputs(2154) <= '0';
    layer0_outputs(2155) <= inputs(85);
    layer0_outputs(2156) <= '0';
    layer0_outputs(2157) <= not(inputs(126));
    layer0_outputs(2158) <= (inputs(74)) xor (inputs(107));
    layer0_outputs(2159) <= (inputs(23)) and not (inputs(142));
    layer0_outputs(2160) <= (inputs(51)) or (inputs(221));
    layer0_outputs(2161) <= (inputs(204)) or (inputs(180));
    layer0_outputs(2162) <= (inputs(232)) and not (inputs(62));
    layer0_outputs(2163) <= (inputs(244)) and not (inputs(134));
    layer0_outputs(2164) <= (inputs(228)) and not (inputs(106));
    layer0_outputs(2165) <= not(inputs(101));
    layer0_outputs(2166) <= not((inputs(62)) or (inputs(79)));
    layer0_outputs(2167) <= not((inputs(211)) or (inputs(203)));
    layer0_outputs(2168) <= not(inputs(50)) or (inputs(0));
    layer0_outputs(2169) <= not((inputs(27)) or (inputs(112)));
    layer0_outputs(2170) <= inputs(82);
    layer0_outputs(2171) <= not(inputs(66));
    layer0_outputs(2172) <= not(inputs(242));
    layer0_outputs(2173) <= not(inputs(202));
    layer0_outputs(2174) <= '1';
    layer0_outputs(2175) <= not(inputs(144));
    layer0_outputs(2176) <= (inputs(156)) or (inputs(130));
    layer0_outputs(2177) <= not((inputs(94)) xor (inputs(8)));
    layer0_outputs(2178) <= not((inputs(1)) xor (inputs(186)));
    layer0_outputs(2179) <= '1';
    layer0_outputs(2180) <= (inputs(92)) and not (inputs(29));
    layer0_outputs(2181) <= inputs(148);
    layer0_outputs(2182) <= not(inputs(64)) or (inputs(199));
    layer0_outputs(2183) <= (inputs(42)) xor (inputs(11));
    layer0_outputs(2184) <= not(inputs(214));
    layer0_outputs(2185) <= (inputs(75)) and (inputs(179));
    layer0_outputs(2186) <= inputs(212);
    layer0_outputs(2187) <= not(inputs(76)) or (inputs(161));
    layer0_outputs(2188) <= inputs(158);
    layer0_outputs(2189) <= (inputs(234)) and not (inputs(5));
    layer0_outputs(2190) <= not((inputs(29)) xor (inputs(115)));
    layer0_outputs(2191) <= (inputs(156)) xor (inputs(221));
    layer0_outputs(2192) <= not(inputs(115)) or (inputs(34));
    layer0_outputs(2193) <= not(inputs(32));
    layer0_outputs(2194) <= inputs(59);
    layer0_outputs(2195) <= (inputs(76)) and not (inputs(71));
    layer0_outputs(2196) <= not((inputs(21)) or (inputs(107)));
    layer0_outputs(2197) <= not(inputs(13)) or (inputs(11));
    layer0_outputs(2198) <= not(inputs(132));
    layer0_outputs(2199) <= not(inputs(197)) or (inputs(182));
    layer0_outputs(2200) <= not(inputs(6));
    layer0_outputs(2201) <= (inputs(254)) xor (inputs(42));
    layer0_outputs(2202) <= not((inputs(163)) or (inputs(229)));
    layer0_outputs(2203) <= not((inputs(187)) or (inputs(45)));
    layer0_outputs(2204) <= not(inputs(181));
    layer0_outputs(2205) <= (inputs(224)) and (inputs(110));
    layer0_outputs(2206) <= (inputs(196)) or (inputs(230));
    layer0_outputs(2207) <= '0';
    layer0_outputs(2208) <= (inputs(73)) and not (inputs(195));
    layer0_outputs(2209) <= inputs(244);
    layer0_outputs(2210) <= (inputs(229)) or (inputs(133));
    layer0_outputs(2211) <= (inputs(28)) or (inputs(151));
    layer0_outputs(2212) <= (inputs(216)) and (inputs(189));
    layer0_outputs(2213) <= not((inputs(139)) or (inputs(189)));
    layer0_outputs(2214) <= not((inputs(85)) or (inputs(246)));
    layer0_outputs(2215) <= (inputs(37)) or (inputs(45));
    layer0_outputs(2216) <= (inputs(239)) and not (inputs(45));
    layer0_outputs(2217) <= not((inputs(177)) or (inputs(33)));
    layer0_outputs(2218) <= not(inputs(131)) or (inputs(248));
    layer0_outputs(2219) <= inputs(146);
    layer0_outputs(2220) <= inputs(206);
    layer0_outputs(2221) <= inputs(128);
    layer0_outputs(2222) <= inputs(25);
    layer0_outputs(2223) <= '1';
    layer0_outputs(2224) <= not((inputs(95)) or (inputs(87)));
    layer0_outputs(2225) <= not((inputs(72)) or (inputs(190)));
    layer0_outputs(2226) <= (inputs(195)) xor (inputs(249));
    layer0_outputs(2227) <= (inputs(24)) and not (inputs(177));
    layer0_outputs(2228) <= inputs(180);
    layer0_outputs(2229) <= not(inputs(4)) or (inputs(254));
    layer0_outputs(2230) <= not(inputs(157));
    layer0_outputs(2231) <= (inputs(9)) xor (inputs(20));
    layer0_outputs(2232) <= not((inputs(191)) or (inputs(167)));
    layer0_outputs(2233) <= not((inputs(86)) or (inputs(54)));
    layer0_outputs(2234) <= '1';
    layer0_outputs(2235) <= not(inputs(145));
    layer0_outputs(2236) <= inputs(185);
    layer0_outputs(2237) <= not((inputs(68)) xor (inputs(80)));
    layer0_outputs(2238) <= not((inputs(80)) xor (inputs(23)));
    layer0_outputs(2239) <= not(inputs(213)) or (inputs(55));
    layer0_outputs(2240) <= not((inputs(148)) and (inputs(230)));
    layer0_outputs(2241) <= inputs(80);
    layer0_outputs(2242) <= (inputs(32)) and (inputs(2));
    layer0_outputs(2243) <= inputs(209);
    layer0_outputs(2244) <= not((inputs(84)) or (inputs(69)));
    layer0_outputs(2245) <= (inputs(56)) and not (inputs(91));
    layer0_outputs(2246) <= not(inputs(166));
    layer0_outputs(2247) <= '1';
    layer0_outputs(2248) <= inputs(200);
    layer0_outputs(2249) <= inputs(239);
    layer0_outputs(2250) <= not((inputs(222)) xor (inputs(103)));
    layer0_outputs(2251) <= not(inputs(203)) or (inputs(238));
    layer0_outputs(2252) <= not(inputs(200));
    layer0_outputs(2253) <= not((inputs(95)) and (inputs(145)));
    layer0_outputs(2254) <= not((inputs(103)) xor (inputs(89)));
    layer0_outputs(2255) <= inputs(90);
    layer0_outputs(2256) <= (inputs(132)) or (inputs(130));
    layer0_outputs(2257) <= not(inputs(170));
    layer0_outputs(2258) <= inputs(10);
    layer0_outputs(2259) <= not((inputs(55)) or (inputs(87)));
    layer0_outputs(2260) <= not((inputs(28)) or (inputs(13)));
    layer0_outputs(2261) <= '1';
    layer0_outputs(2262) <= not(inputs(189));
    layer0_outputs(2263) <= not(inputs(166));
    layer0_outputs(2264) <= (inputs(116)) and not (inputs(216));
    layer0_outputs(2265) <= not((inputs(203)) or (inputs(107)));
    layer0_outputs(2266) <= '1';
    layer0_outputs(2267) <= (inputs(235)) or (inputs(19));
    layer0_outputs(2268) <= (inputs(22)) and not (inputs(1));
    layer0_outputs(2269) <= not((inputs(145)) or (inputs(111)));
    layer0_outputs(2270) <= (inputs(80)) or (inputs(211));
    layer0_outputs(2271) <= not(inputs(19));
    layer0_outputs(2272) <= not((inputs(122)) or (inputs(156)));
    layer0_outputs(2273) <= not(inputs(74));
    layer0_outputs(2274) <= (inputs(159)) and not (inputs(209));
    layer0_outputs(2275) <= (inputs(35)) or (inputs(3));
    layer0_outputs(2276) <= not((inputs(42)) or (inputs(246)));
    layer0_outputs(2277) <= (inputs(65)) or (inputs(208));
    layer0_outputs(2278) <= inputs(88);
    layer0_outputs(2279) <= (inputs(253)) or (inputs(90));
    layer0_outputs(2280) <= (inputs(228)) and not (inputs(74));
    layer0_outputs(2281) <= not(inputs(62));
    layer0_outputs(2282) <= (inputs(57)) or (inputs(21));
    layer0_outputs(2283) <= not(inputs(67));
    layer0_outputs(2284) <= inputs(33);
    layer0_outputs(2285) <= inputs(143);
    layer0_outputs(2286) <= inputs(43);
    layer0_outputs(2287) <= not(inputs(199)) or (inputs(148));
    layer0_outputs(2288) <= not((inputs(188)) and (inputs(222)));
    layer0_outputs(2289) <= not((inputs(118)) or (inputs(133)));
    layer0_outputs(2290) <= not(inputs(252)) or (inputs(96));
    layer0_outputs(2291) <= not(inputs(188));
    layer0_outputs(2292) <= not((inputs(127)) or (inputs(163)));
    layer0_outputs(2293) <= '0';
    layer0_outputs(2294) <= not(inputs(250));
    layer0_outputs(2295) <= inputs(194);
    layer0_outputs(2296) <= (inputs(152)) and (inputs(189));
    layer0_outputs(2297) <= (inputs(17)) or (inputs(20));
    layer0_outputs(2298) <= not(inputs(114)) or (inputs(210));
    layer0_outputs(2299) <= (inputs(92)) or (inputs(98));
    layer0_outputs(2300) <= '0';
    layer0_outputs(2301) <= inputs(40);
    layer0_outputs(2302) <= not(inputs(157));
    layer0_outputs(2303) <= inputs(247);
    layer0_outputs(2304) <= not(inputs(132)) or (inputs(210));
    layer0_outputs(2305) <= not((inputs(240)) or (inputs(89)));
    layer0_outputs(2306) <= (inputs(185)) and not (inputs(30));
    layer0_outputs(2307) <= inputs(245);
    layer0_outputs(2308) <= inputs(183);
    layer0_outputs(2309) <= inputs(98);
    layer0_outputs(2310) <= (inputs(41)) and not (inputs(88));
    layer0_outputs(2311) <= inputs(148);
    layer0_outputs(2312) <= (inputs(145)) xor (inputs(136));
    layer0_outputs(2313) <= not((inputs(218)) or (inputs(238)));
    layer0_outputs(2314) <= inputs(164);
    layer0_outputs(2315) <= inputs(164);
    layer0_outputs(2316) <= (inputs(4)) and not (inputs(232));
    layer0_outputs(2317) <= (inputs(70)) and (inputs(210));
    layer0_outputs(2318) <= '0';
    layer0_outputs(2319) <= (inputs(190)) and not (inputs(191));
    layer0_outputs(2320) <= (inputs(155)) or (inputs(77));
    layer0_outputs(2321) <= inputs(116);
    layer0_outputs(2322) <= not(inputs(130)) or (inputs(197));
    layer0_outputs(2323) <= not(inputs(255));
    layer0_outputs(2324) <= (inputs(236)) xor (inputs(189));
    layer0_outputs(2325) <= not(inputs(84)) or (inputs(222));
    layer0_outputs(2326) <= not(inputs(233));
    layer0_outputs(2327) <= not(inputs(84)) or (inputs(50));
    layer0_outputs(2328) <= inputs(165);
    layer0_outputs(2329) <= (inputs(18)) xor (inputs(155));
    layer0_outputs(2330) <= (inputs(166)) and (inputs(221));
    layer0_outputs(2331) <= not(inputs(162)) or (inputs(31));
    layer0_outputs(2332) <= inputs(237);
    layer0_outputs(2333) <= not(inputs(142));
    layer0_outputs(2334) <= inputs(56);
    layer0_outputs(2335) <= (inputs(51)) and (inputs(106));
    layer0_outputs(2336) <= not((inputs(28)) xor (inputs(59)));
    layer0_outputs(2337) <= (inputs(195)) xor (inputs(5));
    layer0_outputs(2338) <= (inputs(126)) or (inputs(168));
    layer0_outputs(2339) <= (inputs(204)) and not (inputs(20));
    layer0_outputs(2340) <= (inputs(12)) or (inputs(192));
    layer0_outputs(2341) <= (inputs(164)) and not (inputs(192));
    layer0_outputs(2342) <= not(inputs(210));
    layer0_outputs(2343) <= not((inputs(154)) or (inputs(206)));
    layer0_outputs(2344) <= not((inputs(95)) or (inputs(78)));
    layer0_outputs(2345) <= inputs(248);
    layer0_outputs(2346) <= not(inputs(31)) or (inputs(253));
    layer0_outputs(2347) <= inputs(146);
    layer0_outputs(2348) <= (inputs(124)) and not (inputs(222));
    layer0_outputs(2349) <= inputs(134);
    layer0_outputs(2350) <= (inputs(131)) xor (inputs(118));
    layer0_outputs(2351) <= not((inputs(213)) xor (inputs(252)));
    layer0_outputs(2352) <= (inputs(18)) or (inputs(143));
    layer0_outputs(2353) <= not(inputs(107)) or (inputs(8));
    layer0_outputs(2354) <= not((inputs(144)) or (inputs(13)));
    layer0_outputs(2355) <= not(inputs(101));
    layer0_outputs(2356) <= inputs(38);
    layer0_outputs(2357) <= not(inputs(197));
    layer0_outputs(2358) <= not((inputs(188)) and (inputs(72)));
    layer0_outputs(2359) <= (inputs(244)) xor (inputs(126));
    layer0_outputs(2360) <= (inputs(204)) and (inputs(96));
    layer0_outputs(2361) <= (inputs(135)) and not (inputs(209));
    layer0_outputs(2362) <= inputs(181);
    layer0_outputs(2363) <= inputs(184);
    layer0_outputs(2364) <= not(inputs(225)) or (inputs(251));
    layer0_outputs(2365) <= not((inputs(49)) or (inputs(223)));
    layer0_outputs(2366) <= inputs(161);
    layer0_outputs(2367) <= not((inputs(97)) and (inputs(160)));
    layer0_outputs(2368) <= not((inputs(20)) or (inputs(63)));
    layer0_outputs(2369) <= not((inputs(12)) or (inputs(92)));
    layer0_outputs(2370) <= (inputs(41)) or (inputs(126));
    layer0_outputs(2371) <= (inputs(73)) and not (inputs(5));
    layer0_outputs(2372) <= (inputs(157)) or (inputs(145));
    layer0_outputs(2373) <= not((inputs(147)) xor (inputs(171)));
    layer0_outputs(2374) <= not(inputs(115));
    layer0_outputs(2375) <= inputs(90);
    layer0_outputs(2376) <= '1';
    layer0_outputs(2377) <= (inputs(197)) and not (inputs(253));
    layer0_outputs(2378) <= not((inputs(48)) or (inputs(65)));
    layer0_outputs(2379) <= inputs(235);
    layer0_outputs(2380) <= not((inputs(76)) xor (inputs(79)));
    layer0_outputs(2381) <= not((inputs(117)) or (inputs(148)));
    layer0_outputs(2382) <= not(inputs(18));
    layer0_outputs(2383) <= not(inputs(54));
    layer0_outputs(2384) <= not(inputs(194));
    layer0_outputs(2385) <= (inputs(202)) xor (inputs(169));
    layer0_outputs(2386) <= not((inputs(251)) xor (inputs(136)));
    layer0_outputs(2387) <= (inputs(85)) or (inputs(84));
    layer0_outputs(2388) <= inputs(169);
    layer0_outputs(2389) <= inputs(161);
    layer0_outputs(2390) <= not(inputs(243));
    layer0_outputs(2391) <= (inputs(44)) and not (inputs(64));
    layer0_outputs(2392) <= '0';
    layer0_outputs(2393) <= not((inputs(162)) xor (inputs(243)));
    layer0_outputs(2394) <= not(inputs(112));
    layer0_outputs(2395) <= not(inputs(21)) or (inputs(71));
    layer0_outputs(2396) <= inputs(214);
    layer0_outputs(2397) <= not(inputs(31)) or (inputs(217));
    layer0_outputs(2398) <= (inputs(12)) or (inputs(82));
    layer0_outputs(2399) <= '1';
    layer0_outputs(2400) <= not((inputs(39)) or (inputs(138)));
    layer0_outputs(2401) <= inputs(178);
    layer0_outputs(2402) <= inputs(67);
    layer0_outputs(2403) <= not((inputs(248)) or (inputs(193)));
    layer0_outputs(2404) <= not(inputs(126));
    layer0_outputs(2405) <= (inputs(219)) and not (inputs(131));
    layer0_outputs(2406) <= '0';
    layer0_outputs(2407) <= not(inputs(130));
    layer0_outputs(2408) <= not((inputs(105)) or (inputs(7)));
    layer0_outputs(2409) <= (inputs(72)) and not (inputs(192));
    layer0_outputs(2410) <= not(inputs(75));
    layer0_outputs(2411) <= (inputs(9)) and not (inputs(0));
    layer0_outputs(2412) <= inputs(138);
    layer0_outputs(2413) <= not((inputs(91)) xor (inputs(95)));
    layer0_outputs(2414) <= inputs(215);
    layer0_outputs(2415) <= not(inputs(230));
    layer0_outputs(2416) <= not(inputs(222));
    layer0_outputs(2417) <= inputs(67);
    layer0_outputs(2418) <= (inputs(156)) and (inputs(195));
    layer0_outputs(2419) <= not(inputs(76));
    layer0_outputs(2420) <= not(inputs(14));
    layer0_outputs(2421) <= not((inputs(194)) or (inputs(179)));
    layer0_outputs(2422) <= inputs(116);
    layer0_outputs(2423) <= (inputs(112)) and not (inputs(192));
    layer0_outputs(2424) <= (inputs(132)) and not (inputs(225));
    layer0_outputs(2425) <= (inputs(131)) or (inputs(163));
    layer0_outputs(2426) <= not(inputs(206)) or (inputs(114));
    layer0_outputs(2427) <= (inputs(112)) and not (inputs(49));
    layer0_outputs(2428) <= not((inputs(36)) xor (inputs(20)));
    layer0_outputs(2429) <= (inputs(19)) or (inputs(122));
    layer0_outputs(2430) <= inputs(7);
    layer0_outputs(2431) <= '0';
    layer0_outputs(2432) <= not(inputs(159)) or (inputs(165));
    layer0_outputs(2433) <= inputs(82);
    layer0_outputs(2434) <= not((inputs(85)) xor (inputs(127)));
    layer0_outputs(2435) <= inputs(214);
    layer0_outputs(2436) <= '0';
    layer0_outputs(2437) <= (inputs(73)) or (inputs(47));
    layer0_outputs(2438) <= not((inputs(20)) xor (inputs(94)));
    layer0_outputs(2439) <= (inputs(166)) and not (inputs(46));
    layer0_outputs(2440) <= inputs(9);
    layer0_outputs(2441) <= (inputs(14)) or (inputs(208));
    layer0_outputs(2442) <= (inputs(172)) or (inputs(237));
    layer0_outputs(2443) <= (inputs(178)) and not (inputs(95));
    layer0_outputs(2444) <= not(inputs(91)) or (inputs(216));
    layer0_outputs(2445) <= not(inputs(101));
    layer0_outputs(2446) <= (inputs(19)) and not (inputs(229));
    layer0_outputs(2447) <= (inputs(247)) and not (inputs(253));
    layer0_outputs(2448) <= not(inputs(56));
    layer0_outputs(2449) <= not(inputs(254));
    layer0_outputs(2450) <= (inputs(240)) xor (inputs(152));
    layer0_outputs(2451) <= (inputs(78)) and not (inputs(18));
    layer0_outputs(2452) <= (inputs(252)) or (inputs(102));
    layer0_outputs(2453) <= (inputs(36)) or (inputs(45));
    layer0_outputs(2454) <= (inputs(130)) xor (inputs(53));
    layer0_outputs(2455) <= not((inputs(70)) or (inputs(16)));
    layer0_outputs(2456) <= (inputs(89)) xor (inputs(169));
    layer0_outputs(2457) <= (inputs(100)) or (inputs(124));
    layer0_outputs(2458) <= not(inputs(182)) or (inputs(90));
    layer0_outputs(2459) <= not(inputs(117)) or (inputs(246));
    layer0_outputs(2460) <= (inputs(35)) xor (inputs(125));
    layer0_outputs(2461) <= (inputs(122)) and not (inputs(16));
    layer0_outputs(2462) <= inputs(139);
    layer0_outputs(2463) <= (inputs(255)) or (inputs(89));
    layer0_outputs(2464) <= (inputs(126)) and (inputs(243));
    layer0_outputs(2465) <= not(inputs(246));
    layer0_outputs(2466) <= not((inputs(153)) xor (inputs(214)));
    layer0_outputs(2467) <= (inputs(195)) and not (inputs(251));
    layer0_outputs(2468) <= (inputs(231)) or (inputs(118));
    layer0_outputs(2469) <= not((inputs(237)) and (inputs(74)));
    layer0_outputs(2470) <= not((inputs(64)) xor (inputs(188)));
    layer0_outputs(2471) <= not((inputs(48)) xor (inputs(8)));
    layer0_outputs(2472) <= not((inputs(103)) or (inputs(213)));
    layer0_outputs(2473) <= not(inputs(40));
    layer0_outputs(2474) <= not(inputs(188));
    layer0_outputs(2475) <= not(inputs(57));
    layer0_outputs(2476) <= not(inputs(187));
    layer0_outputs(2477) <= not((inputs(229)) or (inputs(219)));
    layer0_outputs(2478) <= (inputs(25)) and not (inputs(116));
    layer0_outputs(2479) <= '0';
    layer0_outputs(2480) <= (inputs(223)) or (inputs(205));
    layer0_outputs(2481) <= (inputs(19)) xor (inputs(81));
    layer0_outputs(2482) <= (inputs(84)) and not (inputs(224));
    layer0_outputs(2483) <= '0';
    layer0_outputs(2484) <= inputs(122);
    layer0_outputs(2485) <= inputs(29);
    layer0_outputs(2486) <= not((inputs(110)) xor (inputs(90)));
    layer0_outputs(2487) <= inputs(93);
    layer0_outputs(2488) <= not(inputs(21));
    layer0_outputs(2489) <= inputs(147);
    layer0_outputs(2490) <= inputs(212);
    layer0_outputs(2491) <= '1';
    layer0_outputs(2492) <= (inputs(49)) xor (inputs(21));
    layer0_outputs(2493) <= inputs(133);
    layer0_outputs(2494) <= not(inputs(129)) or (inputs(136));
    layer0_outputs(2495) <= inputs(123);
    layer0_outputs(2496) <= (inputs(117)) and not (inputs(12));
    layer0_outputs(2497) <= inputs(55);
    layer0_outputs(2498) <= (inputs(6)) and not (inputs(172));
    layer0_outputs(2499) <= (inputs(144)) xor (inputs(249));
    layer0_outputs(2500) <= not(inputs(179)) or (inputs(89));
    layer0_outputs(2501) <= inputs(137);
    layer0_outputs(2502) <= not((inputs(1)) or (inputs(156)));
    layer0_outputs(2503) <= not((inputs(122)) or (inputs(28)));
    layer0_outputs(2504) <= not(inputs(26)) or (inputs(212));
    layer0_outputs(2505) <= not((inputs(166)) or (inputs(147)));
    layer0_outputs(2506) <= not(inputs(10)) or (inputs(0));
    layer0_outputs(2507) <= not(inputs(183));
    layer0_outputs(2508) <= not((inputs(133)) xor (inputs(20)));
    layer0_outputs(2509) <= not((inputs(144)) xor (inputs(210)));
    layer0_outputs(2510) <= not((inputs(126)) xor (inputs(144)));
    layer0_outputs(2511) <= not(inputs(227));
    layer0_outputs(2512) <= not((inputs(76)) or (inputs(224)));
    layer0_outputs(2513) <= '1';
    layer0_outputs(2514) <= (inputs(76)) and not (inputs(128));
    layer0_outputs(2515) <= inputs(68);
    layer0_outputs(2516) <= inputs(233);
    layer0_outputs(2517) <= not(inputs(237)) or (inputs(74));
    layer0_outputs(2518) <= not(inputs(196));
    layer0_outputs(2519) <= '1';
    layer0_outputs(2520) <= not((inputs(35)) or (inputs(167)));
    layer0_outputs(2521) <= not(inputs(140));
    layer0_outputs(2522) <= (inputs(54)) or (inputs(220));
    layer0_outputs(2523) <= not(inputs(227)) or (inputs(18));
    layer0_outputs(2524) <= not(inputs(169));
    layer0_outputs(2525) <= not(inputs(187));
    layer0_outputs(2526) <= (inputs(67)) xor (inputs(151));
    layer0_outputs(2527) <= (inputs(200)) or (inputs(111));
    layer0_outputs(2528) <= (inputs(246)) or (inputs(40));
    layer0_outputs(2529) <= not((inputs(70)) and (inputs(245)));
    layer0_outputs(2530) <= not((inputs(45)) or (inputs(109)));
    layer0_outputs(2531) <= not(inputs(236));
    layer0_outputs(2532) <= (inputs(34)) and not (inputs(6));
    layer0_outputs(2533) <= not((inputs(184)) or (inputs(159)));
    layer0_outputs(2534) <= not(inputs(242)) or (inputs(220));
    layer0_outputs(2535) <= not(inputs(87));
    layer0_outputs(2536) <= inputs(198);
    layer0_outputs(2537) <= not((inputs(216)) or (inputs(224)));
    layer0_outputs(2538) <= not(inputs(122));
    layer0_outputs(2539) <= not(inputs(131));
    layer0_outputs(2540) <= not(inputs(94)) or (inputs(20));
    layer0_outputs(2541) <= (inputs(67)) and not (inputs(175));
    layer0_outputs(2542) <= not((inputs(156)) or (inputs(157)));
    layer0_outputs(2543) <= not((inputs(155)) or (inputs(31)));
    layer0_outputs(2544) <= '1';
    layer0_outputs(2545) <= inputs(55);
    layer0_outputs(2546) <= not((inputs(89)) or (inputs(66)));
    layer0_outputs(2547) <= not(inputs(177));
    layer0_outputs(2548) <= not(inputs(45)) or (inputs(167));
    layer0_outputs(2549) <= (inputs(26)) and not (inputs(183));
    layer0_outputs(2550) <= (inputs(199)) and not (inputs(28));
    layer0_outputs(2551) <= not((inputs(245)) and (inputs(179)));
    layer0_outputs(2552) <= not(inputs(66));
    layer0_outputs(2553) <= (inputs(129)) or (inputs(42));
    layer0_outputs(2554) <= not((inputs(221)) or (inputs(213)));
    layer0_outputs(2555) <= inputs(86);
    layer0_outputs(2556) <= inputs(37);
    layer0_outputs(2557) <= not(inputs(70));
    layer0_outputs(2558) <= not(inputs(115)) or (inputs(222));
    layer0_outputs(2559) <= not(inputs(130));
    layer0_outputs(2560) <= not(inputs(100)) or (inputs(48));
    layer0_outputs(2561) <= not((inputs(9)) or (inputs(43)));
    layer0_outputs(2562) <= inputs(189);
    layer0_outputs(2563) <= (inputs(135)) and not (inputs(140));
    layer0_outputs(2564) <= inputs(44);
    layer0_outputs(2565) <= (inputs(76)) and (inputs(90));
    layer0_outputs(2566) <= not((inputs(212)) or (inputs(32)));
    layer0_outputs(2567) <= not((inputs(186)) and (inputs(113)));
    layer0_outputs(2568) <= not(inputs(214));
    layer0_outputs(2569) <= not((inputs(69)) or (inputs(129)));
    layer0_outputs(2570) <= (inputs(213)) or (inputs(205));
    layer0_outputs(2571) <= inputs(160);
    layer0_outputs(2572) <= (inputs(97)) xor (inputs(86));
    layer0_outputs(2573) <= (inputs(233)) and not (inputs(93));
    layer0_outputs(2574) <= not(inputs(37));
    layer0_outputs(2575) <= (inputs(37)) and (inputs(255));
    layer0_outputs(2576) <= not(inputs(226)) or (inputs(140));
    layer0_outputs(2577) <= not(inputs(92)) or (inputs(126));
    layer0_outputs(2578) <= not(inputs(162));
    layer0_outputs(2579) <= (inputs(242)) xor (inputs(143));
    layer0_outputs(2580) <= '0';
    layer0_outputs(2581) <= not(inputs(109)) or (inputs(232));
    layer0_outputs(2582) <= not(inputs(255)) or (inputs(49));
    layer0_outputs(2583) <= '1';
    layer0_outputs(2584) <= not(inputs(45));
    layer0_outputs(2585) <= not((inputs(47)) and (inputs(118)));
    layer0_outputs(2586) <= inputs(170);
    layer0_outputs(2587) <= inputs(74);
    layer0_outputs(2588) <= (inputs(129)) and not (inputs(253));
    layer0_outputs(2589) <= not((inputs(85)) and (inputs(75)));
    layer0_outputs(2590) <= (inputs(223)) or (inputs(208));
    layer0_outputs(2591) <= not(inputs(95));
    layer0_outputs(2592) <= (inputs(55)) and not (inputs(103));
    layer0_outputs(2593) <= inputs(147);
    layer0_outputs(2594) <= not(inputs(203));
    layer0_outputs(2595) <= (inputs(127)) xor (inputs(52));
    layer0_outputs(2596) <= not(inputs(41));
    layer0_outputs(2597) <= not(inputs(212)) or (inputs(50));
    layer0_outputs(2598) <= not(inputs(177));
    layer0_outputs(2599) <= not((inputs(148)) and (inputs(236)));
    layer0_outputs(2600) <= not((inputs(145)) or (inputs(166)));
    layer0_outputs(2601) <= inputs(38);
    layer0_outputs(2602) <= not((inputs(35)) or (inputs(88)));
    layer0_outputs(2603) <= not(inputs(116)) or (inputs(225));
    layer0_outputs(2604) <= (inputs(27)) and (inputs(15));
    layer0_outputs(2605) <= (inputs(92)) and not (inputs(26));
    layer0_outputs(2606) <= not(inputs(228));
    layer0_outputs(2607) <= (inputs(114)) or (inputs(99));
    layer0_outputs(2608) <= inputs(151);
    layer0_outputs(2609) <= inputs(244);
    layer0_outputs(2610) <= inputs(46);
    layer0_outputs(2611) <= not((inputs(19)) xor (inputs(254)));
    layer0_outputs(2612) <= not(inputs(174));
    layer0_outputs(2613) <= inputs(78);
    layer0_outputs(2614) <= inputs(71);
    layer0_outputs(2615) <= not(inputs(175));
    layer0_outputs(2616) <= not(inputs(99));
    layer0_outputs(2617) <= '0';
    layer0_outputs(2618) <= not(inputs(118));
    layer0_outputs(2619) <= not(inputs(8)) or (inputs(199));
    layer0_outputs(2620) <= inputs(228);
    layer0_outputs(2621) <= not((inputs(210)) or (inputs(164)));
    layer0_outputs(2622) <= '0';
    layer0_outputs(2623) <= inputs(152);
    layer0_outputs(2624) <= inputs(233);
    layer0_outputs(2625) <= not(inputs(32)) or (inputs(8));
    layer0_outputs(2626) <= inputs(220);
    layer0_outputs(2627) <= not((inputs(22)) xor (inputs(73)));
    layer0_outputs(2628) <= inputs(52);
    layer0_outputs(2629) <= not((inputs(158)) and (inputs(114)));
    layer0_outputs(2630) <= (inputs(27)) xor (inputs(5));
    layer0_outputs(2631) <= (inputs(133)) and not (inputs(10));
    layer0_outputs(2632) <= not((inputs(243)) xor (inputs(227)));
    layer0_outputs(2633) <= (inputs(250)) and not (inputs(64));
    layer0_outputs(2634) <= inputs(37);
    layer0_outputs(2635) <= inputs(9);
    layer0_outputs(2636) <= (inputs(253)) or (inputs(166));
    layer0_outputs(2637) <= (inputs(103)) and (inputs(132));
    layer0_outputs(2638) <= (inputs(137)) and not (inputs(239));
    layer0_outputs(2639) <= not((inputs(117)) xor (inputs(161)));
    layer0_outputs(2640) <= (inputs(119)) and not (inputs(127));
    layer0_outputs(2641) <= inputs(229);
    layer0_outputs(2642) <= (inputs(78)) and not (inputs(239));
    layer0_outputs(2643) <= not((inputs(47)) and (inputs(145)));
    layer0_outputs(2644) <= not(inputs(54)) or (inputs(28));
    layer0_outputs(2645) <= '1';
    layer0_outputs(2646) <= '1';
    layer0_outputs(2647) <= (inputs(184)) and not (inputs(87));
    layer0_outputs(2648) <= not(inputs(62)) or (inputs(253));
    layer0_outputs(2649) <= (inputs(221)) xor (inputs(60));
    layer0_outputs(2650) <= (inputs(209)) xor (inputs(181));
    layer0_outputs(2651) <= not((inputs(167)) xor (inputs(140)));
    layer0_outputs(2652) <= inputs(189);
    layer0_outputs(2653) <= not(inputs(97));
    layer0_outputs(2654) <= '0';
    layer0_outputs(2655) <= (inputs(242)) or (inputs(171));
    layer0_outputs(2656) <= inputs(183);
    layer0_outputs(2657) <= not((inputs(155)) or (inputs(185)));
    layer0_outputs(2658) <= not(inputs(88));
    layer0_outputs(2659) <= not(inputs(190));
    layer0_outputs(2660) <= (inputs(101)) and not (inputs(4));
    layer0_outputs(2661) <= not(inputs(17));
    layer0_outputs(2662) <= not(inputs(75)) or (inputs(200));
    layer0_outputs(2663) <= not(inputs(16)) or (inputs(124));
    layer0_outputs(2664) <= not((inputs(202)) or (inputs(132)));
    layer0_outputs(2665) <= not(inputs(82));
    layer0_outputs(2666) <= not((inputs(40)) and (inputs(22)));
    layer0_outputs(2667) <= not(inputs(91));
    layer0_outputs(2668) <= (inputs(73)) and not (inputs(177));
    layer0_outputs(2669) <= inputs(113);
    layer0_outputs(2670) <= (inputs(121)) xor (inputs(88));
    layer0_outputs(2671) <= not((inputs(146)) or (inputs(178)));
    layer0_outputs(2672) <= not(inputs(225));
    layer0_outputs(2673) <= not(inputs(122));
    layer0_outputs(2674) <= (inputs(210)) and not (inputs(42));
    layer0_outputs(2675) <= (inputs(254)) or (inputs(131));
    layer0_outputs(2676) <= not((inputs(56)) xor (inputs(43)));
    layer0_outputs(2677) <= inputs(4);
    layer0_outputs(2678) <= not((inputs(127)) xor (inputs(108)));
    layer0_outputs(2679) <= (inputs(181)) xor (inputs(138));
    layer0_outputs(2680) <= inputs(2);
    layer0_outputs(2681) <= not((inputs(231)) or (inputs(128)));
    layer0_outputs(2682) <= (inputs(164)) and not (inputs(128));
    layer0_outputs(2683) <= not(inputs(147)) or (inputs(0));
    layer0_outputs(2684) <= not(inputs(195)) or (inputs(115));
    layer0_outputs(2685) <= '0';
    layer0_outputs(2686) <= not((inputs(23)) and (inputs(27)));
    layer0_outputs(2687) <= '0';
    layer0_outputs(2688) <= not(inputs(190));
    layer0_outputs(2689) <= (inputs(154)) and (inputs(147));
    layer0_outputs(2690) <= (inputs(77)) xor (inputs(57));
    layer0_outputs(2691) <= '1';
    layer0_outputs(2692) <= not((inputs(192)) and (inputs(102)));
    layer0_outputs(2693) <= not((inputs(241)) or (inputs(189)));
    layer0_outputs(2694) <= '0';
    layer0_outputs(2695) <= not((inputs(243)) or (inputs(51)));
    layer0_outputs(2696) <= not(inputs(86));
    layer0_outputs(2697) <= not((inputs(246)) xor (inputs(19)));
    layer0_outputs(2698) <= inputs(10);
    layer0_outputs(2699) <= (inputs(163)) and not (inputs(60));
    layer0_outputs(2700) <= not(inputs(69)) or (inputs(178));
    layer0_outputs(2701) <= not(inputs(61));
    layer0_outputs(2702) <= inputs(161);
    layer0_outputs(2703) <= not(inputs(60));
    layer0_outputs(2704) <= not(inputs(21));
    layer0_outputs(2705) <= '0';
    layer0_outputs(2706) <= inputs(102);
    layer0_outputs(2707) <= not((inputs(188)) or (inputs(54)));
    layer0_outputs(2708) <= (inputs(133)) and (inputs(91));
    layer0_outputs(2709) <= not(inputs(167)) or (inputs(52));
    layer0_outputs(2710) <= inputs(249);
    layer0_outputs(2711) <= (inputs(162)) xor (inputs(158));
    layer0_outputs(2712) <= not(inputs(10));
    layer0_outputs(2713) <= not(inputs(206));
    layer0_outputs(2714) <= not(inputs(219));
    layer0_outputs(2715) <= inputs(166);
    layer0_outputs(2716) <= not((inputs(219)) or (inputs(84)));
    layer0_outputs(2717) <= not((inputs(178)) and (inputs(73)));
    layer0_outputs(2718) <= not(inputs(102));
    layer0_outputs(2719) <= not(inputs(146));
    layer0_outputs(2720) <= (inputs(17)) or (inputs(101));
    layer0_outputs(2721) <= not((inputs(74)) or (inputs(7)));
    layer0_outputs(2722) <= (inputs(20)) and not (inputs(200));
    layer0_outputs(2723) <= not((inputs(40)) xor (inputs(176)));
    layer0_outputs(2724) <= (inputs(123)) and (inputs(176));
    layer0_outputs(2725) <= (inputs(20)) or (inputs(115));
    layer0_outputs(2726) <= inputs(172);
    layer0_outputs(2727) <= (inputs(71)) and not (inputs(241));
    layer0_outputs(2728) <= (inputs(142)) and not (inputs(252));
    layer0_outputs(2729) <= (inputs(239)) xor (inputs(136));
    layer0_outputs(2730) <= not((inputs(139)) or (inputs(138)));
    layer0_outputs(2731) <= (inputs(131)) xor (inputs(50));
    layer0_outputs(2732) <= not((inputs(248)) xor (inputs(204)));
    layer0_outputs(2733) <= not((inputs(31)) or (inputs(241)));
    layer0_outputs(2734) <= (inputs(12)) or (inputs(17));
    layer0_outputs(2735) <= inputs(87);
    layer0_outputs(2736) <= (inputs(250)) and (inputs(249));
    layer0_outputs(2737) <= not((inputs(67)) and (inputs(64)));
    layer0_outputs(2738) <= '0';
    layer0_outputs(2739) <= not(inputs(39));
    layer0_outputs(2740) <= not((inputs(11)) and (inputs(240)));
    layer0_outputs(2741) <= (inputs(28)) xor (inputs(45));
    layer0_outputs(2742) <= not(inputs(227));
    layer0_outputs(2743) <= not((inputs(149)) or (inputs(196)));
    layer0_outputs(2744) <= inputs(105);
    layer0_outputs(2745) <= not(inputs(137));
    layer0_outputs(2746) <= '1';
    layer0_outputs(2747) <= not(inputs(154));
    layer0_outputs(2748) <= (inputs(170)) and (inputs(138));
    layer0_outputs(2749) <= not(inputs(83));
    layer0_outputs(2750) <= not(inputs(24)) or (inputs(174));
    layer0_outputs(2751) <= (inputs(24)) and not (inputs(151));
    layer0_outputs(2752) <= (inputs(221)) xor (inputs(210));
    layer0_outputs(2753) <= not((inputs(195)) or (inputs(8)));
    layer0_outputs(2754) <= not(inputs(232)) or (inputs(118));
    layer0_outputs(2755) <= not(inputs(99));
    layer0_outputs(2756) <= not(inputs(109));
    layer0_outputs(2757) <= (inputs(15)) or (inputs(103));
    layer0_outputs(2758) <= inputs(91);
    layer0_outputs(2759) <= not(inputs(228));
    layer0_outputs(2760) <= not(inputs(60));
    layer0_outputs(2761) <= (inputs(140)) and not (inputs(15));
    layer0_outputs(2762) <= '1';
    layer0_outputs(2763) <= inputs(210);
    layer0_outputs(2764) <= inputs(180);
    layer0_outputs(2765) <= not((inputs(97)) xor (inputs(87)));
    layer0_outputs(2766) <= not(inputs(88)) or (inputs(16));
    layer0_outputs(2767) <= (inputs(104)) or (inputs(99));
    layer0_outputs(2768) <= not(inputs(111)) or (inputs(242));
    layer0_outputs(2769) <= not(inputs(236)) or (inputs(14));
    layer0_outputs(2770) <= not((inputs(224)) or (inputs(187)));
    layer0_outputs(2771) <= (inputs(25)) xor (inputs(73));
    layer0_outputs(2772) <= not(inputs(0)) or (inputs(118));
    layer0_outputs(2773) <= (inputs(223)) and not (inputs(80));
    layer0_outputs(2774) <= not(inputs(106));
    layer0_outputs(2775) <= (inputs(144)) and not (inputs(94));
    layer0_outputs(2776) <= not(inputs(140)) or (inputs(223));
    layer0_outputs(2777) <= not(inputs(162));
    layer0_outputs(2778) <= inputs(122);
    layer0_outputs(2779) <= not(inputs(209));
    layer0_outputs(2780) <= inputs(145);
    layer0_outputs(2781) <= (inputs(199)) or (inputs(174));
    layer0_outputs(2782) <= not((inputs(130)) or (inputs(245)));
    layer0_outputs(2783) <= not((inputs(253)) or (inputs(88)));
    layer0_outputs(2784) <= (inputs(174)) xor (inputs(156));
    layer0_outputs(2785) <= not((inputs(71)) or (inputs(255)));
    layer0_outputs(2786) <= not((inputs(233)) or (inputs(213)));
    layer0_outputs(2787) <= not((inputs(243)) or (inputs(197)));
    layer0_outputs(2788) <= '1';
    layer0_outputs(2789) <= not(inputs(22));
    layer0_outputs(2790) <= not((inputs(20)) xor (inputs(37)));
    layer0_outputs(2791) <= inputs(153);
    layer0_outputs(2792) <= (inputs(140)) or (inputs(69));
    layer0_outputs(2793) <= not(inputs(224));
    layer0_outputs(2794) <= (inputs(42)) and not (inputs(123));
    layer0_outputs(2795) <= (inputs(9)) xor (inputs(72));
    layer0_outputs(2796) <= not((inputs(168)) and (inputs(214)));
    layer0_outputs(2797) <= not(inputs(31));
    layer0_outputs(2798) <= not((inputs(149)) xor (inputs(63)));
    layer0_outputs(2799) <= (inputs(24)) and not (inputs(190));
    layer0_outputs(2800) <= not(inputs(151));
    layer0_outputs(2801) <= not(inputs(106));
    layer0_outputs(2802) <= (inputs(101)) xor (inputs(11));
    layer0_outputs(2803) <= not((inputs(126)) or (inputs(143)));
    layer0_outputs(2804) <= not(inputs(53));
    layer0_outputs(2805) <= not((inputs(71)) and (inputs(192)));
    layer0_outputs(2806) <= not(inputs(18));
    layer0_outputs(2807) <= (inputs(6)) and not (inputs(251));
    layer0_outputs(2808) <= (inputs(223)) and not (inputs(234));
    layer0_outputs(2809) <= not((inputs(116)) and (inputs(80)));
    layer0_outputs(2810) <= inputs(173);
    layer0_outputs(2811) <= not((inputs(88)) or (inputs(163)));
    layer0_outputs(2812) <= not((inputs(38)) or (inputs(170)));
    layer0_outputs(2813) <= inputs(59);
    layer0_outputs(2814) <= (inputs(12)) or (inputs(0));
    layer0_outputs(2815) <= not(inputs(161));
    layer0_outputs(2816) <= inputs(211);
    layer0_outputs(2817) <= inputs(164);
    layer0_outputs(2818) <= not(inputs(84));
    layer0_outputs(2819) <= (inputs(155)) and not (inputs(94));
    layer0_outputs(2820) <= not((inputs(27)) xor (inputs(142)));
    layer0_outputs(2821) <= not(inputs(89)) or (inputs(232));
    layer0_outputs(2822) <= not(inputs(120)) or (inputs(174));
    layer0_outputs(2823) <= (inputs(36)) or (inputs(173));
    layer0_outputs(2824) <= not(inputs(141));
    layer0_outputs(2825) <= inputs(170);
    layer0_outputs(2826) <= inputs(76);
    layer0_outputs(2827) <= inputs(167);
    layer0_outputs(2828) <= (inputs(161)) or (inputs(199));
    layer0_outputs(2829) <= not(inputs(217));
    layer0_outputs(2830) <= '0';
    layer0_outputs(2831) <= not(inputs(123));
    layer0_outputs(2832) <= inputs(61);
    layer0_outputs(2833) <= (inputs(194)) and not (inputs(205));
    layer0_outputs(2834) <= (inputs(40)) or (inputs(157));
    layer0_outputs(2835) <= (inputs(204)) and not (inputs(60));
    layer0_outputs(2836) <= inputs(96);
    layer0_outputs(2837) <= (inputs(158)) and (inputs(142));
    layer0_outputs(2838) <= inputs(154);
    layer0_outputs(2839) <= not(inputs(44)) or (inputs(38));
    layer0_outputs(2840) <= not((inputs(252)) xor (inputs(155)));
    layer0_outputs(2841) <= (inputs(218)) and not (inputs(240));
    layer0_outputs(2842) <= not(inputs(40));
    layer0_outputs(2843) <= not(inputs(242)) or (inputs(151));
    layer0_outputs(2844) <= not(inputs(132));
    layer0_outputs(2845) <= not(inputs(114));
    layer0_outputs(2846) <= inputs(111);
    layer0_outputs(2847) <= not(inputs(121));
    layer0_outputs(2848) <= inputs(217);
    layer0_outputs(2849) <= (inputs(168)) or (inputs(133));
    layer0_outputs(2850) <= inputs(153);
    layer0_outputs(2851) <= inputs(161);
    layer0_outputs(2852) <= (inputs(171)) xor (inputs(203));
    layer0_outputs(2853) <= (inputs(74)) and not (inputs(1));
    layer0_outputs(2854) <= (inputs(107)) and not (inputs(80));
    layer0_outputs(2855) <= inputs(198);
    layer0_outputs(2856) <= not((inputs(250)) xor (inputs(187)));
    layer0_outputs(2857) <= (inputs(132)) and (inputs(38));
    layer0_outputs(2858) <= not(inputs(141));
    layer0_outputs(2859) <= not(inputs(177)) or (inputs(214));
    layer0_outputs(2860) <= not((inputs(202)) or (inputs(227)));
    layer0_outputs(2861) <= not(inputs(71));
    layer0_outputs(2862) <= (inputs(9)) and not (inputs(185));
    layer0_outputs(2863) <= inputs(113);
    layer0_outputs(2864) <= not(inputs(232)) or (inputs(15));
    layer0_outputs(2865) <= not(inputs(178));
    layer0_outputs(2866) <= not((inputs(243)) or (inputs(36)));
    layer0_outputs(2867) <= '1';
    layer0_outputs(2868) <= not(inputs(165));
    layer0_outputs(2869) <= (inputs(227)) and (inputs(134));
    layer0_outputs(2870) <= not(inputs(145)) or (inputs(135));
    layer0_outputs(2871) <= not((inputs(156)) xor (inputs(106)));
    layer0_outputs(2872) <= (inputs(212)) and not (inputs(253));
    layer0_outputs(2873) <= (inputs(244)) and not (inputs(128));
    layer0_outputs(2874) <= (inputs(233)) and not (inputs(240));
    layer0_outputs(2875) <= not(inputs(122)) or (inputs(32));
    layer0_outputs(2876) <= inputs(211);
    layer0_outputs(2877) <= not((inputs(132)) xor (inputs(69)));
    layer0_outputs(2878) <= (inputs(52)) xor (inputs(104));
    layer0_outputs(2879) <= (inputs(140)) or (inputs(150));
    layer0_outputs(2880) <= not(inputs(122));
    layer0_outputs(2881) <= (inputs(197)) and not (inputs(32));
    layer0_outputs(2882) <= not(inputs(192));
    layer0_outputs(2883) <= not((inputs(254)) and (inputs(127)));
    layer0_outputs(2884) <= (inputs(68)) and not (inputs(165));
    layer0_outputs(2885) <= '0';
    layer0_outputs(2886) <= (inputs(95)) xor (inputs(245));
    layer0_outputs(2887) <= (inputs(90)) xor (inputs(2));
    layer0_outputs(2888) <= not(inputs(168)) or (inputs(159));
    layer0_outputs(2889) <= inputs(122);
    layer0_outputs(2890) <= (inputs(47)) or (inputs(215));
    layer0_outputs(2891) <= inputs(182);
    layer0_outputs(2892) <= (inputs(88)) and not (inputs(66));
    layer0_outputs(2893) <= not(inputs(61));
    layer0_outputs(2894) <= '1';
    layer0_outputs(2895) <= (inputs(148)) and not (inputs(33));
    layer0_outputs(2896) <= not(inputs(141));
    layer0_outputs(2897) <= not((inputs(237)) or (inputs(235)));
    layer0_outputs(2898) <= not((inputs(234)) xor (inputs(195)));
    layer0_outputs(2899) <= not((inputs(150)) or (inputs(81)));
    layer0_outputs(2900) <= not(inputs(134)) or (inputs(187));
    layer0_outputs(2901) <= not((inputs(71)) or (inputs(235)));
    layer0_outputs(2902) <= (inputs(133)) or (inputs(121));
    layer0_outputs(2903) <= (inputs(91)) and (inputs(175));
    layer0_outputs(2904) <= inputs(16);
    layer0_outputs(2905) <= (inputs(203)) xor (inputs(18));
    layer0_outputs(2906) <= (inputs(103)) or (inputs(46));
    layer0_outputs(2907) <= not(inputs(177)) or (inputs(128));
    layer0_outputs(2908) <= not((inputs(108)) or (inputs(208)));
    layer0_outputs(2909) <= not((inputs(16)) or (inputs(26)));
    layer0_outputs(2910) <= not(inputs(2));
    layer0_outputs(2911) <= not(inputs(160));
    layer0_outputs(2912) <= inputs(125);
    layer0_outputs(2913) <= not((inputs(7)) xor (inputs(195)));
    layer0_outputs(2914) <= not(inputs(197)) or (inputs(32));
    layer0_outputs(2915) <= (inputs(121)) and not (inputs(113));
    layer0_outputs(2916) <= not(inputs(144)) or (inputs(128));
    layer0_outputs(2917) <= not((inputs(170)) or (inputs(179)));
    layer0_outputs(2918) <= not((inputs(10)) xor (inputs(143)));
    layer0_outputs(2919) <= not(inputs(239));
    layer0_outputs(2920) <= inputs(149);
    layer0_outputs(2921) <= (inputs(133)) or (inputs(187));
    layer0_outputs(2922) <= (inputs(228)) and not (inputs(90));
    layer0_outputs(2923) <= not(inputs(40));
    layer0_outputs(2924) <= not(inputs(107)) or (inputs(206));
    layer0_outputs(2925) <= (inputs(149)) or (inputs(134));
    layer0_outputs(2926) <= (inputs(128)) or (inputs(132));
    layer0_outputs(2927) <= not(inputs(182));
    layer0_outputs(2928) <= (inputs(223)) and not (inputs(143));
    layer0_outputs(2929) <= not(inputs(219));
    layer0_outputs(2930) <= inputs(192);
    layer0_outputs(2931) <= not((inputs(245)) or (inputs(215)));
    layer0_outputs(2932) <= not(inputs(178));
    layer0_outputs(2933) <= '1';
    layer0_outputs(2934) <= not(inputs(140));
    layer0_outputs(2935) <= not((inputs(21)) or (inputs(2)));
    layer0_outputs(2936) <= not(inputs(114));
    layer0_outputs(2937) <= not((inputs(239)) or (inputs(147)));
    layer0_outputs(2938) <= (inputs(100)) and not (inputs(55));
    layer0_outputs(2939) <= not(inputs(122));
    layer0_outputs(2940) <= not(inputs(22));
    layer0_outputs(2941) <= (inputs(22)) or (inputs(124));
    layer0_outputs(2942) <= not(inputs(110));
    layer0_outputs(2943) <= not(inputs(150));
    layer0_outputs(2944) <= not(inputs(206)) or (inputs(179));
    layer0_outputs(2945) <= not(inputs(227));
    layer0_outputs(2946) <= not((inputs(90)) xor (inputs(43)));
    layer0_outputs(2947) <= not(inputs(183)) or (inputs(5));
    layer0_outputs(2948) <= inputs(204);
    layer0_outputs(2949) <= not(inputs(194));
    layer0_outputs(2950) <= (inputs(62)) and not (inputs(165));
    layer0_outputs(2951) <= not(inputs(182)) or (inputs(186));
    layer0_outputs(2952) <= not(inputs(11));
    layer0_outputs(2953) <= inputs(149);
    layer0_outputs(2954) <= not(inputs(250));
    layer0_outputs(2955) <= not(inputs(180));
    layer0_outputs(2956) <= not(inputs(242));
    layer0_outputs(2957) <= not(inputs(191)) or (inputs(123));
    layer0_outputs(2958) <= not(inputs(142));
    layer0_outputs(2959) <= not(inputs(253)) or (inputs(197));
    layer0_outputs(2960) <= not(inputs(212));
    layer0_outputs(2961) <= not(inputs(142)) or (inputs(240));
    layer0_outputs(2962) <= not((inputs(147)) or (inputs(237)));
    layer0_outputs(2963) <= (inputs(127)) or (inputs(236));
    layer0_outputs(2964) <= (inputs(233)) xor (inputs(144));
    layer0_outputs(2965) <= not((inputs(10)) or (inputs(80)));
    layer0_outputs(2966) <= not((inputs(92)) or (inputs(207)));
    layer0_outputs(2967) <= not((inputs(75)) or (inputs(253)));
    layer0_outputs(2968) <= not(inputs(85));
    layer0_outputs(2969) <= not((inputs(89)) xor (inputs(189)));
    layer0_outputs(2970) <= not((inputs(34)) or (inputs(153)));
    layer0_outputs(2971) <= not((inputs(246)) or (inputs(74)));
    layer0_outputs(2972) <= not(inputs(172)) or (inputs(66));
    layer0_outputs(2973) <= '1';
    layer0_outputs(2974) <= not((inputs(144)) and (inputs(162)));
    layer0_outputs(2975) <= inputs(62);
    layer0_outputs(2976) <= inputs(83);
    layer0_outputs(2977) <= inputs(180);
    layer0_outputs(2978) <= not(inputs(247)) or (inputs(255));
    layer0_outputs(2979) <= inputs(182);
    layer0_outputs(2980) <= not((inputs(61)) or (inputs(103)));
    layer0_outputs(2981) <= not((inputs(65)) and (inputs(247)));
    layer0_outputs(2982) <= (inputs(29)) or (inputs(221));
    layer0_outputs(2983) <= not(inputs(132)) or (inputs(214));
    layer0_outputs(2984) <= not((inputs(171)) or (inputs(180)));
    layer0_outputs(2985) <= inputs(125);
    layer0_outputs(2986) <= inputs(225);
    layer0_outputs(2987) <= not((inputs(138)) or (inputs(192)));
    layer0_outputs(2988) <= inputs(70);
    layer0_outputs(2989) <= not((inputs(155)) or (inputs(114)));
    layer0_outputs(2990) <= not(inputs(12));
    layer0_outputs(2991) <= (inputs(128)) and not (inputs(147));
    layer0_outputs(2992) <= not((inputs(28)) xor (inputs(103)));
    layer0_outputs(2993) <= (inputs(205)) and not (inputs(159));
    layer0_outputs(2994) <= (inputs(72)) and not (inputs(35));
    layer0_outputs(2995) <= not((inputs(82)) xor (inputs(25)));
    layer0_outputs(2996) <= not(inputs(39));
    layer0_outputs(2997) <= (inputs(0)) and not (inputs(199));
    layer0_outputs(2998) <= (inputs(78)) and not (inputs(3));
    layer0_outputs(2999) <= not(inputs(23));
    layer0_outputs(3000) <= not((inputs(28)) or (inputs(84)));
    layer0_outputs(3001) <= not((inputs(148)) and (inputs(75)));
    layer0_outputs(3002) <= not((inputs(234)) or (inputs(96)));
    layer0_outputs(3003) <= not(inputs(166));
    layer0_outputs(3004) <= not((inputs(179)) or (inputs(97)));
    layer0_outputs(3005) <= not(inputs(99));
    layer0_outputs(3006) <= (inputs(57)) and not (inputs(21));
    layer0_outputs(3007) <= (inputs(26)) and not (inputs(132));
    layer0_outputs(3008) <= '0';
    layer0_outputs(3009) <= not(inputs(90));
    layer0_outputs(3010) <= inputs(121);
    layer0_outputs(3011) <= inputs(15);
    layer0_outputs(3012) <= inputs(148);
    layer0_outputs(3013) <= (inputs(53)) and not (inputs(238));
    layer0_outputs(3014) <= '0';
    layer0_outputs(3015) <= not((inputs(89)) xor (inputs(13)));
    layer0_outputs(3016) <= '0';
    layer0_outputs(3017) <= inputs(106);
    layer0_outputs(3018) <= inputs(158);
    layer0_outputs(3019) <= '1';
    layer0_outputs(3020) <= not((inputs(81)) and (inputs(20)));
    layer0_outputs(3021) <= not((inputs(70)) xor (inputs(87)));
    layer0_outputs(3022) <= inputs(79);
    layer0_outputs(3023) <= (inputs(90)) or (inputs(109));
    layer0_outputs(3024) <= (inputs(73)) xor (inputs(208));
    layer0_outputs(3025) <= not((inputs(128)) and (inputs(44)));
    layer0_outputs(3026) <= (inputs(223)) or (inputs(229));
    layer0_outputs(3027) <= (inputs(88)) or (inputs(103));
    layer0_outputs(3028) <= (inputs(175)) and not (inputs(204));
    layer0_outputs(3029) <= (inputs(34)) and not (inputs(184));
    layer0_outputs(3030) <= not(inputs(247));
    layer0_outputs(3031) <= inputs(75);
    layer0_outputs(3032) <= (inputs(5)) xor (inputs(187));
    layer0_outputs(3033) <= (inputs(55)) xor (inputs(123));
    layer0_outputs(3034) <= not((inputs(75)) and (inputs(121)));
    layer0_outputs(3035) <= not((inputs(77)) or (inputs(205)));
    layer0_outputs(3036) <= (inputs(66)) and not (inputs(197));
    layer0_outputs(3037) <= not(inputs(99)) or (inputs(32));
    layer0_outputs(3038) <= not(inputs(19));
    layer0_outputs(3039) <= (inputs(127)) or (inputs(42));
    layer0_outputs(3040) <= (inputs(242)) and (inputs(222));
    layer0_outputs(3041) <= inputs(211);
    layer0_outputs(3042) <= not(inputs(149)) or (inputs(240));
    layer0_outputs(3043) <= inputs(249);
    layer0_outputs(3044) <= not((inputs(146)) and (inputs(130)));
    layer0_outputs(3045) <= (inputs(152)) and not (inputs(159));
    layer0_outputs(3046) <= (inputs(43)) and not (inputs(210));
    layer0_outputs(3047) <= (inputs(154)) or (inputs(101));
    layer0_outputs(3048) <= (inputs(96)) and not (inputs(159));
    layer0_outputs(3049) <= not((inputs(56)) and (inputs(77)));
    layer0_outputs(3050) <= (inputs(16)) xor (inputs(58));
    layer0_outputs(3051) <= not((inputs(0)) and (inputs(1)));
    layer0_outputs(3052) <= inputs(192);
    layer0_outputs(3053) <= not(inputs(72));
    layer0_outputs(3054) <= not(inputs(17));
    layer0_outputs(3055) <= not((inputs(149)) and (inputs(178)));
    layer0_outputs(3056) <= inputs(229);
    layer0_outputs(3057) <= (inputs(153)) and not (inputs(32));
    layer0_outputs(3058) <= (inputs(112)) or (inputs(130));
    layer0_outputs(3059) <= inputs(107);
    layer0_outputs(3060) <= not(inputs(242));
    layer0_outputs(3061) <= not((inputs(121)) xor (inputs(195)));
    layer0_outputs(3062) <= inputs(220);
    layer0_outputs(3063) <= (inputs(149)) or (inputs(148));
    layer0_outputs(3064) <= (inputs(6)) or (inputs(126));
    layer0_outputs(3065) <= (inputs(118)) and not (inputs(16));
    layer0_outputs(3066) <= inputs(161);
    layer0_outputs(3067) <= inputs(200);
    layer0_outputs(3068) <= '0';
    layer0_outputs(3069) <= (inputs(160)) and not (inputs(115));
    layer0_outputs(3070) <= not(inputs(101));
    layer0_outputs(3071) <= '0';
    layer0_outputs(3072) <= not(inputs(120)) or (inputs(155));
    layer0_outputs(3073) <= not((inputs(39)) and (inputs(127)));
    layer0_outputs(3074) <= inputs(84);
    layer0_outputs(3075) <= (inputs(201)) and not (inputs(14));
    layer0_outputs(3076) <= '1';
    layer0_outputs(3077) <= not(inputs(147));
    layer0_outputs(3078) <= inputs(150);
    layer0_outputs(3079) <= not((inputs(65)) or (inputs(72)));
    layer0_outputs(3080) <= not(inputs(123));
    layer0_outputs(3081) <= not((inputs(156)) xor (inputs(185)));
    layer0_outputs(3082) <= (inputs(127)) xor (inputs(189));
    layer0_outputs(3083) <= not((inputs(142)) or (inputs(245)));
    layer0_outputs(3084) <= inputs(131);
    layer0_outputs(3085) <= not(inputs(129));
    layer0_outputs(3086) <= not(inputs(212));
    layer0_outputs(3087) <= (inputs(87)) xor (inputs(140));
    layer0_outputs(3088) <= inputs(210);
    layer0_outputs(3089) <= not(inputs(193)) or (inputs(203));
    layer0_outputs(3090) <= not(inputs(163));
    layer0_outputs(3091) <= (inputs(242)) xor (inputs(165));
    layer0_outputs(3092) <= not(inputs(98));
    layer0_outputs(3093) <= '1';
    layer0_outputs(3094) <= inputs(73);
    layer0_outputs(3095) <= not(inputs(243));
    layer0_outputs(3096) <= not(inputs(28));
    layer0_outputs(3097) <= (inputs(98)) and not (inputs(13));
    layer0_outputs(3098) <= inputs(22);
    layer0_outputs(3099) <= inputs(86);
    layer0_outputs(3100) <= (inputs(134)) xor (inputs(89));
    layer0_outputs(3101) <= not(inputs(215)) or (inputs(128));
    layer0_outputs(3102) <= (inputs(217)) or (inputs(111));
    layer0_outputs(3103) <= not(inputs(227));
    layer0_outputs(3104) <= '1';
    layer0_outputs(3105) <= not(inputs(64));
    layer0_outputs(3106) <= not((inputs(20)) or (inputs(67)));
    layer0_outputs(3107) <= (inputs(142)) or (inputs(96));
    layer0_outputs(3108) <= (inputs(26)) and not (inputs(171));
    layer0_outputs(3109) <= inputs(191);
    layer0_outputs(3110) <= not(inputs(230));
    layer0_outputs(3111) <= inputs(9);
    layer0_outputs(3112) <= not(inputs(163));
    layer0_outputs(3113) <= not(inputs(230)) or (inputs(169));
    layer0_outputs(3114) <= '0';
    layer0_outputs(3115) <= (inputs(175)) and not (inputs(89));
    layer0_outputs(3116) <= not((inputs(73)) xor (inputs(11)));
    layer0_outputs(3117) <= (inputs(197)) xor (inputs(149));
    layer0_outputs(3118) <= not(inputs(197)) or (inputs(36));
    layer0_outputs(3119) <= not(inputs(132)) or (inputs(254));
    layer0_outputs(3120) <= '0';
    layer0_outputs(3121) <= not(inputs(139));
    layer0_outputs(3122) <= (inputs(22)) xor (inputs(13));
    layer0_outputs(3123) <= inputs(25);
    layer0_outputs(3124) <= not(inputs(169));
    layer0_outputs(3125) <= (inputs(87)) or (inputs(215));
    layer0_outputs(3126) <= (inputs(10)) xor (inputs(250));
    layer0_outputs(3127) <= (inputs(51)) and not (inputs(159));
    layer0_outputs(3128) <= '1';
    layer0_outputs(3129) <= not((inputs(8)) or (inputs(171)));
    layer0_outputs(3130) <= inputs(79);
    layer0_outputs(3131) <= (inputs(121)) and not (inputs(64));
    layer0_outputs(3132) <= (inputs(186)) and not (inputs(123));
    layer0_outputs(3133) <= (inputs(109)) or (inputs(110));
    layer0_outputs(3134) <= not(inputs(188)) or (inputs(241));
    layer0_outputs(3135) <= not(inputs(42)) or (inputs(172));
    layer0_outputs(3136) <= not((inputs(232)) xor (inputs(241)));
    layer0_outputs(3137) <= inputs(146);
    layer0_outputs(3138) <= not(inputs(25));
    layer0_outputs(3139) <= not((inputs(189)) or (inputs(71)));
    layer0_outputs(3140) <= not((inputs(66)) and (inputs(59)));
    layer0_outputs(3141) <= inputs(215);
    layer0_outputs(3142) <= (inputs(5)) and not (inputs(96));
    layer0_outputs(3143) <= (inputs(228)) and not (inputs(235));
    layer0_outputs(3144) <= not((inputs(221)) xor (inputs(174)));
    layer0_outputs(3145) <= not(inputs(129)) or (inputs(253));
    layer0_outputs(3146) <= not(inputs(108)) or (inputs(213));
    layer0_outputs(3147) <= not(inputs(217)) or (inputs(153));
    layer0_outputs(3148) <= (inputs(100)) and (inputs(238));
    layer0_outputs(3149) <= not((inputs(65)) or (inputs(34)));
    layer0_outputs(3150) <= inputs(6);
    layer0_outputs(3151) <= not(inputs(115)) or (inputs(33));
    layer0_outputs(3152) <= (inputs(64)) xor (inputs(12));
    layer0_outputs(3153) <= (inputs(34)) or (inputs(154));
    layer0_outputs(3154) <= not((inputs(139)) or (inputs(108)));
    layer0_outputs(3155) <= (inputs(225)) and not (inputs(12));
    layer0_outputs(3156) <= (inputs(69)) or (inputs(124));
    layer0_outputs(3157) <= (inputs(36)) and (inputs(43));
    layer0_outputs(3158) <= inputs(193);
    layer0_outputs(3159) <= inputs(152);
    layer0_outputs(3160) <= not(inputs(222));
    layer0_outputs(3161) <= (inputs(169)) and not (inputs(128));
    layer0_outputs(3162) <= (inputs(174)) and (inputs(52));
    layer0_outputs(3163) <= not((inputs(3)) or (inputs(185)));
    layer0_outputs(3164) <= not(inputs(68));
    layer0_outputs(3165) <= not(inputs(92)) or (inputs(172));
    layer0_outputs(3166) <= not((inputs(193)) or (inputs(167)));
    layer0_outputs(3167) <= (inputs(149)) or (inputs(177));
    layer0_outputs(3168) <= inputs(103);
    layer0_outputs(3169) <= not(inputs(72)) or (inputs(47));
    layer0_outputs(3170) <= not(inputs(147));
    layer0_outputs(3171) <= not(inputs(252));
    layer0_outputs(3172) <= not(inputs(36));
    layer0_outputs(3173) <= not(inputs(79));
    layer0_outputs(3174) <= '0';
    layer0_outputs(3175) <= not(inputs(52));
    layer0_outputs(3176) <= not((inputs(134)) xor (inputs(154)));
    layer0_outputs(3177) <= not(inputs(177));
    layer0_outputs(3178) <= (inputs(64)) or (inputs(184));
    layer0_outputs(3179) <= (inputs(58)) and not (inputs(240));
    layer0_outputs(3180) <= (inputs(177)) xor (inputs(167));
    layer0_outputs(3181) <= (inputs(109)) xor (inputs(78));
    layer0_outputs(3182) <= not(inputs(132));
    layer0_outputs(3183) <= inputs(137);
    layer0_outputs(3184) <= not(inputs(182)) or (inputs(110));
    layer0_outputs(3185) <= not(inputs(225));
    layer0_outputs(3186) <= (inputs(213)) or (inputs(28));
    layer0_outputs(3187) <= not(inputs(121)) or (inputs(24));
    layer0_outputs(3188) <= (inputs(22)) xor (inputs(173));
    layer0_outputs(3189) <= not((inputs(141)) and (inputs(99)));
    layer0_outputs(3190) <= not((inputs(25)) and (inputs(104)));
    layer0_outputs(3191) <= (inputs(117)) or (inputs(224));
    layer0_outputs(3192) <= not((inputs(57)) and (inputs(117)));
    layer0_outputs(3193) <= (inputs(170)) and not (inputs(26));
    layer0_outputs(3194) <= inputs(29);
    layer0_outputs(3195) <= inputs(89);
    layer0_outputs(3196) <= not((inputs(148)) or (inputs(172)));
    layer0_outputs(3197) <= not((inputs(175)) xor (inputs(96)));
    layer0_outputs(3198) <= (inputs(228)) and not (inputs(102));
    layer0_outputs(3199) <= not((inputs(16)) or (inputs(196)));
    layer0_outputs(3200) <= not((inputs(108)) xor (inputs(43)));
    layer0_outputs(3201) <= inputs(193);
    layer0_outputs(3202) <= (inputs(222)) and not (inputs(113));
    layer0_outputs(3203) <= inputs(235);
    layer0_outputs(3204) <= not(inputs(13)) or (inputs(91));
    layer0_outputs(3205) <= inputs(89);
    layer0_outputs(3206) <= not((inputs(198)) or (inputs(75)));
    layer0_outputs(3207) <= not((inputs(243)) or (inputs(192)));
    layer0_outputs(3208) <= (inputs(187)) or (inputs(234));
    layer0_outputs(3209) <= inputs(204);
    layer0_outputs(3210) <= '1';
    layer0_outputs(3211) <= not((inputs(184)) xor (inputs(173)));
    layer0_outputs(3212) <= not((inputs(234)) and (inputs(10)));
    layer0_outputs(3213) <= not((inputs(188)) or (inputs(96)));
    layer0_outputs(3214) <= not(inputs(127));
    layer0_outputs(3215) <= inputs(7);
    layer0_outputs(3216) <= '0';
    layer0_outputs(3217) <= not(inputs(59));
    layer0_outputs(3218) <= (inputs(169)) and not (inputs(97));
    layer0_outputs(3219) <= (inputs(235)) or (inputs(111));
    layer0_outputs(3220) <= not((inputs(212)) or (inputs(212)));
    layer0_outputs(3221) <= not((inputs(115)) or (inputs(138)));
    layer0_outputs(3222) <= not((inputs(80)) or (inputs(50)));
    layer0_outputs(3223) <= not((inputs(169)) or (inputs(15)));
    layer0_outputs(3224) <= not((inputs(42)) or (inputs(232)));
    layer0_outputs(3225) <= inputs(101);
    layer0_outputs(3226) <= not((inputs(76)) and (inputs(43)));
    layer0_outputs(3227) <= not(inputs(147));
    layer0_outputs(3228) <= not((inputs(142)) or (inputs(70)));
    layer0_outputs(3229) <= (inputs(130)) and not (inputs(102));
    layer0_outputs(3230) <= inputs(23);
    layer0_outputs(3231) <= (inputs(54)) or (inputs(160));
    layer0_outputs(3232) <= (inputs(231)) or (inputs(241));
    layer0_outputs(3233) <= not(inputs(70));
    layer0_outputs(3234) <= not(inputs(185)) or (inputs(125));
    layer0_outputs(3235) <= inputs(155);
    layer0_outputs(3236) <= (inputs(185)) or (inputs(236));
    layer0_outputs(3237) <= (inputs(92)) and not (inputs(149));
    layer0_outputs(3238) <= not(inputs(107)) or (inputs(135));
    layer0_outputs(3239) <= not((inputs(240)) xor (inputs(171)));
    layer0_outputs(3240) <= not((inputs(35)) xor (inputs(12)));
    layer0_outputs(3241) <= (inputs(159)) or (inputs(22));
    layer0_outputs(3242) <= (inputs(28)) and not (inputs(42));
    layer0_outputs(3243) <= not(inputs(135));
    layer0_outputs(3244) <= (inputs(250)) and (inputs(231));
    layer0_outputs(3245) <= not(inputs(94));
    layer0_outputs(3246) <= not((inputs(188)) and (inputs(46)));
    layer0_outputs(3247) <= (inputs(85)) and not (inputs(173));
    layer0_outputs(3248) <= not((inputs(117)) xor (inputs(128)));
    layer0_outputs(3249) <= (inputs(120)) or (inputs(129));
    layer0_outputs(3250) <= (inputs(180)) xor (inputs(8));
    layer0_outputs(3251) <= not(inputs(149));
    layer0_outputs(3252) <= not(inputs(7)) or (inputs(159));
    layer0_outputs(3253) <= not(inputs(64)) or (inputs(113));
    layer0_outputs(3254) <= not((inputs(141)) or (inputs(250)));
    layer0_outputs(3255) <= (inputs(234)) and not (inputs(137));
    layer0_outputs(3256) <= not((inputs(151)) or (inputs(178)));
    layer0_outputs(3257) <= inputs(175);
    layer0_outputs(3258) <= not((inputs(205)) or (inputs(103)));
    layer0_outputs(3259) <= not(inputs(54));
    layer0_outputs(3260) <= not((inputs(106)) or (inputs(120)));
    layer0_outputs(3261) <= inputs(71);
    layer0_outputs(3262) <= not((inputs(149)) xor (inputs(145)));
    layer0_outputs(3263) <= not(inputs(30)) or (inputs(237));
    layer0_outputs(3264) <= (inputs(235)) and not (inputs(50));
    layer0_outputs(3265) <= (inputs(197)) and not (inputs(43));
    layer0_outputs(3266) <= not(inputs(94));
    layer0_outputs(3267) <= (inputs(42)) xor (inputs(232));
    layer0_outputs(3268) <= (inputs(241)) or (inputs(137));
    layer0_outputs(3269) <= (inputs(178)) or (inputs(219));
    layer0_outputs(3270) <= not((inputs(247)) or (inputs(132)));
    layer0_outputs(3271) <= not((inputs(16)) xor (inputs(108)));
    layer0_outputs(3272) <= (inputs(99)) and not (inputs(136));
    layer0_outputs(3273) <= not((inputs(35)) xor (inputs(129)));
    layer0_outputs(3274) <= not(inputs(184)) or (inputs(11));
    layer0_outputs(3275) <= not((inputs(168)) xor (inputs(147)));
    layer0_outputs(3276) <= not(inputs(21)) or (inputs(174));
    layer0_outputs(3277) <= not((inputs(229)) or (inputs(227)));
    layer0_outputs(3278) <= (inputs(41)) or (inputs(30));
    layer0_outputs(3279) <= (inputs(240)) or (inputs(198));
    layer0_outputs(3280) <= inputs(107);
    layer0_outputs(3281) <= not(inputs(116));
    layer0_outputs(3282) <= (inputs(202)) or (inputs(85));
    layer0_outputs(3283) <= not((inputs(169)) xor (inputs(252)));
    layer0_outputs(3284) <= (inputs(192)) xor (inputs(83));
    layer0_outputs(3285) <= not((inputs(100)) xor (inputs(237)));
    layer0_outputs(3286) <= not(inputs(61));
    layer0_outputs(3287) <= (inputs(186)) and not (inputs(19));
    layer0_outputs(3288) <= not((inputs(241)) xor (inputs(214)));
    layer0_outputs(3289) <= not((inputs(231)) xor (inputs(111)));
    layer0_outputs(3290) <= (inputs(138)) xor (inputs(144));
    layer0_outputs(3291) <= inputs(163);
    layer0_outputs(3292) <= not((inputs(255)) or (inputs(147)));
    layer0_outputs(3293) <= not(inputs(194)) or (inputs(158));
    layer0_outputs(3294) <= not(inputs(152)) or (inputs(52));
    layer0_outputs(3295) <= inputs(172);
    layer0_outputs(3296) <= (inputs(144)) or (inputs(65));
    layer0_outputs(3297) <= not(inputs(93)) or (inputs(134));
    layer0_outputs(3298) <= (inputs(203)) and not (inputs(15));
    layer0_outputs(3299) <= not(inputs(77)) or (inputs(240));
    layer0_outputs(3300) <= not(inputs(90));
    layer0_outputs(3301) <= (inputs(109)) or (inputs(150));
    layer0_outputs(3302) <= (inputs(153)) and not (inputs(213));
    layer0_outputs(3303) <= (inputs(66)) and not (inputs(127));
    layer0_outputs(3304) <= (inputs(137)) or (inputs(237));
    layer0_outputs(3305) <= (inputs(214)) or (inputs(236));
    layer0_outputs(3306) <= (inputs(146)) and (inputs(241));
    layer0_outputs(3307) <= not(inputs(70));
    layer0_outputs(3308) <= (inputs(180)) xor (inputs(83));
    layer0_outputs(3309) <= inputs(98);
    layer0_outputs(3310) <= (inputs(131)) and (inputs(200));
    layer0_outputs(3311) <= not(inputs(190));
    layer0_outputs(3312) <= inputs(95);
    layer0_outputs(3313) <= not(inputs(193));
    layer0_outputs(3314) <= (inputs(96)) and not (inputs(10));
    layer0_outputs(3315) <= not(inputs(115));
    layer0_outputs(3316) <= not(inputs(248));
    layer0_outputs(3317) <= inputs(21);
    layer0_outputs(3318) <= not((inputs(218)) and (inputs(218)));
    layer0_outputs(3319) <= not((inputs(164)) and (inputs(201)));
    layer0_outputs(3320) <= (inputs(178)) and not (inputs(255));
    layer0_outputs(3321) <= not(inputs(240));
    layer0_outputs(3322) <= not((inputs(145)) xor (inputs(133)));
    layer0_outputs(3323) <= not((inputs(146)) or (inputs(164)));
    layer0_outputs(3324) <= not(inputs(9));
    layer0_outputs(3325) <= (inputs(178)) or (inputs(220));
    layer0_outputs(3326) <= (inputs(3)) xor (inputs(16));
    layer0_outputs(3327) <= not((inputs(239)) or (inputs(112)));
    layer0_outputs(3328) <= not(inputs(141)) or (inputs(191));
    layer0_outputs(3329) <= not(inputs(1)) or (inputs(254));
    layer0_outputs(3330) <= not((inputs(235)) xor (inputs(221)));
    layer0_outputs(3331) <= (inputs(35)) or (inputs(178));
    layer0_outputs(3332) <= not(inputs(198));
    layer0_outputs(3333) <= (inputs(197)) and not (inputs(66));
    layer0_outputs(3334) <= not((inputs(83)) xor (inputs(70)));
    layer0_outputs(3335) <= not(inputs(229));
    layer0_outputs(3336) <= inputs(106);
    layer0_outputs(3337) <= inputs(157);
    layer0_outputs(3338) <= not(inputs(185)) or (inputs(152));
    layer0_outputs(3339) <= (inputs(0)) xor (inputs(138));
    layer0_outputs(3340) <= (inputs(147)) or (inputs(129));
    layer0_outputs(3341) <= not(inputs(70));
    layer0_outputs(3342) <= not(inputs(13)) or (inputs(57));
    layer0_outputs(3343) <= (inputs(148)) xor (inputs(29));
    layer0_outputs(3344) <= (inputs(124)) or (inputs(203));
    layer0_outputs(3345) <= '1';
    layer0_outputs(3346) <= (inputs(104)) xor (inputs(90));
    layer0_outputs(3347) <= not(inputs(253)) or (inputs(86));
    layer0_outputs(3348) <= not((inputs(49)) xor (inputs(4)));
    layer0_outputs(3349) <= not((inputs(222)) or (inputs(235)));
    layer0_outputs(3350) <= not((inputs(76)) or (inputs(65)));
    layer0_outputs(3351) <= not(inputs(17));
    layer0_outputs(3352) <= inputs(178);
    layer0_outputs(3353) <= not(inputs(42));
    layer0_outputs(3354) <= '1';
    layer0_outputs(3355) <= not(inputs(213));
    layer0_outputs(3356) <= (inputs(180)) and not (inputs(211));
    layer0_outputs(3357) <= (inputs(66)) or (inputs(16));
    layer0_outputs(3358) <= not(inputs(117));
    layer0_outputs(3359) <= inputs(200);
    layer0_outputs(3360) <= not(inputs(213)) or (inputs(73));
    layer0_outputs(3361) <= not((inputs(27)) or (inputs(18)));
    layer0_outputs(3362) <= not((inputs(147)) xor (inputs(38)));
    layer0_outputs(3363) <= not((inputs(57)) xor (inputs(22)));
    layer0_outputs(3364) <= (inputs(222)) and not (inputs(66));
    layer0_outputs(3365) <= inputs(212);
    layer0_outputs(3366) <= not(inputs(80));
    layer0_outputs(3367) <= (inputs(79)) and not (inputs(243));
    layer0_outputs(3368) <= inputs(176);
    layer0_outputs(3369) <= not(inputs(5));
    layer0_outputs(3370) <= inputs(252);
    layer0_outputs(3371) <= not((inputs(158)) or (inputs(96)));
    layer0_outputs(3372) <= not(inputs(153));
    layer0_outputs(3373) <= inputs(206);
    layer0_outputs(3374) <= (inputs(20)) xor (inputs(186));
    layer0_outputs(3375) <= inputs(182);
    layer0_outputs(3376) <= not(inputs(216));
    layer0_outputs(3377) <= (inputs(178)) xor (inputs(195));
    layer0_outputs(3378) <= inputs(139);
    layer0_outputs(3379) <= not(inputs(128));
    layer0_outputs(3380) <= not((inputs(59)) xor (inputs(135)));
    layer0_outputs(3381) <= (inputs(109)) and not (inputs(80));
    layer0_outputs(3382) <= inputs(68);
    layer0_outputs(3383) <= not(inputs(180));
    layer0_outputs(3384) <= (inputs(240)) xor (inputs(152));
    layer0_outputs(3385) <= (inputs(33)) or (inputs(105));
    layer0_outputs(3386) <= (inputs(249)) and (inputs(30));
    layer0_outputs(3387) <= not(inputs(66)) or (inputs(48));
    layer0_outputs(3388) <= (inputs(68)) or (inputs(12));
    layer0_outputs(3389) <= not(inputs(224));
    layer0_outputs(3390) <= not(inputs(155));
    layer0_outputs(3391) <= (inputs(91)) or (inputs(99));
    layer0_outputs(3392) <= (inputs(146)) and not (inputs(135));
    layer0_outputs(3393) <= not((inputs(16)) or (inputs(62)));
    layer0_outputs(3394) <= not(inputs(81)) or (inputs(219));
    layer0_outputs(3395) <= not((inputs(90)) or (inputs(152)));
    layer0_outputs(3396) <= '1';
    layer0_outputs(3397) <= not((inputs(158)) or (inputs(176)));
    layer0_outputs(3398) <= not((inputs(47)) or (inputs(83)));
    layer0_outputs(3399) <= not(inputs(232));
    layer0_outputs(3400) <= '0';
    layer0_outputs(3401) <= (inputs(60)) or (inputs(77));
    layer0_outputs(3402) <= (inputs(193)) and not (inputs(31));
    layer0_outputs(3403) <= not(inputs(11));
    layer0_outputs(3404) <= inputs(40);
    layer0_outputs(3405) <= not(inputs(14));
    layer0_outputs(3406) <= (inputs(176)) or (inputs(26));
    layer0_outputs(3407) <= (inputs(210)) and not (inputs(96));
    layer0_outputs(3408) <= not((inputs(20)) or (inputs(209)));
    layer0_outputs(3409) <= not(inputs(112));
    layer0_outputs(3410) <= inputs(101);
    layer0_outputs(3411) <= (inputs(228)) and not (inputs(161));
    layer0_outputs(3412) <= not(inputs(247));
    layer0_outputs(3413) <= not(inputs(164));
    layer0_outputs(3414) <= (inputs(233)) and not (inputs(13));
    layer0_outputs(3415) <= inputs(95);
    layer0_outputs(3416) <= not(inputs(74)) or (inputs(14));
    layer0_outputs(3417) <= inputs(89);
    layer0_outputs(3418) <= not((inputs(133)) or (inputs(206)));
    layer0_outputs(3419) <= not((inputs(35)) xor (inputs(3)));
    layer0_outputs(3420) <= (inputs(91)) and not (inputs(225));
    layer0_outputs(3421) <= not(inputs(164));
    layer0_outputs(3422) <= (inputs(38)) xor (inputs(10));
    layer0_outputs(3423) <= inputs(157);
    layer0_outputs(3424) <= (inputs(147)) xor (inputs(81));
    layer0_outputs(3425) <= not((inputs(69)) xor (inputs(21)));
    layer0_outputs(3426) <= not((inputs(128)) xor (inputs(92)));
    layer0_outputs(3427) <= (inputs(123)) and not (inputs(88));
    layer0_outputs(3428) <= '0';
    layer0_outputs(3429) <= not(inputs(4));
    layer0_outputs(3430) <= not(inputs(187));
    layer0_outputs(3431) <= not((inputs(130)) or (inputs(239)));
    layer0_outputs(3432) <= (inputs(120)) and not (inputs(125));
    layer0_outputs(3433) <= not(inputs(69)) or (inputs(93));
    layer0_outputs(3434) <= (inputs(42)) and not (inputs(236));
    layer0_outputs(3435) <= not(inputs(220)) or (inputs(46));
    layer0_outputs(3436) <= not(inputs(140));
    layer0_outputs(3437) <= (inputs(8)) and not (inputs(26));
    layer0_outputs(3438) <= not(inputs(38)) or (inputs(237));
    layer0_outputs(3439) <= not((inputs(0)) or (inputs(19)));
    layer0_outputs(3440) <= (inputs(4)) and not (inputs(221));
    layer0_outputs(3441) <= (inputs(9)) and not (inputs(134));
    layer0_outputs(3442) <= (inputs(50)) and not (inputs(255));
    layer0_outputs(3443) <= '1';
    layer0_outputs(3444) <= not((inputs(175)) or (inputs(36)));
    layer0_outputs(3445) <= not(inputs(133)) or (inputs(0));
    layer0_outputs(3446) <= not(inputs(105)) or (inputs(191));
    layer0_outputs(3447) <= not(inputs(115)) or (inputs(255));
    layer0_outputs(3448) <= (inputs(206)) or (inputs(185));
    layer0_outputs(3449) <= (inputs(74)) or (inputs(106));
    layer0_outputs(3450) <= (inputs(217)) and not (inputs(138));
    layer0_outputs(3451) <= not(inputs(8));
    layer0_outputs(3452) <= inputs(83);
    layer0_outputs(3453) <= not(inputs(58)) or (inputs(194));
    layer0_outputs(3454) <= (inputs(202)) and not (inputs(139));
    layer0_outputs(3455) <= inputs(165);
    layer0_outputs(3456) <= not((inputs(110)) or (inputs(135)));
    layer0_outputs(3457) <= (inputs(160)) xor (inputs(183));
    layer0_outputs(3458) <= inputs(107);
    layer0_outputs(3459) <= not((inputs(110)) or (inputs(147)));
    layer0_outputs(3460) <= (inputs(235)) and not (inputs(143));
    layer0_outputs(3461) <= (inputs(137)) and not (inputs(129));
    layer0_outputs(3462) <= not((inputs(52)) or (inputs(31)));
    layer0_outputs(3463) <= (inputs(76)) and not (inputs(242));
    layer0_outputs(3464) <= not(inputs(144));
    layer0_outputs(3465) <= not((inputs(0)) or (inputs(141)));
    layer0_outputs(3466) <= not(inputs(8)) or (inputs(135));
    layer0_outputs(3467) <= not(inputs(13)) or (inputs(207));
    layer0_outputs(3468) <= inputs(154);
    layer0_outputs(3469) <= not(inputs(235)) or (inputs(118));
    layer0_outputs(3470) <= inputs(194);
    layer0_outputs(3471) <= not(inputs(14)) or (inputs(38));
    layer0_outputs(3472) <= not(inputs(232));
    layer0_outputs(3473) <= (inputs(107)) and not (inputs(103));
    layer0_outputs(3474) <= not((inputs(182)) xor (inputs(139)));
    layer0_outputs(3475) <= not((inputs(65)) or (inputs(253)));
    layer0_outputs(3476) <= (inputs(21)) or (inputs(27));
    layer0_outputs(3477) <= not(inputs(2));
    layer0_outputs(3478) <= (inputs(122)) and not (inputs(56));
    layer0_outputs(3479) <= inputs(77);
    layer0_outputs(3480) <= (inputs(72)) and not (inputs(2));
    layer0_outputs(3481) <= not(inputs(217)) or (inputs(39));
    layer0_outputs(3482) <= not((inputs(79)) or (inputs(63)));
    layer0_outputs(3483) <= (inputs(110)) and not (inputs(189));
    layer0_outputs(3484) <= (inputs(243)) or (inputs(141));
    layer0_outputs(3485) <= inputs(99);
    layer0_outputs(3486) <= inputs(154);
    layer0_outputs(3487) <= (inputs(71)) and (inputs(72));
    layer0_outputs(3488) <= inputs(140);
    layer0_outputs(3489) <= not(inputs(158)) or (inputs(43));
    layer0_outputs(3490) <= not(inputs(122)) or (inputs(73));
    layer0_outputs(3491) <= (inputs(67)) or (inputs(130));
    layer0_outputs(3492) <= (inputs(148)) and not (inputs(58));
    layer0_outputs(3493) <= not(inputs(252));
    layer0_outputs(3494) <= not(inputs(217));
    layer0_outputs(3495) <= not(inputs(225)) or (inputs(30));
    layer0_outputs(3496) <= inputs(86);
    layer0_outputs(3497) <= not((inputs(80)) xor (inputs(170)));
    layer0_outputs(3498) <= not((inputs(180)) or (inputs(171)));
    layer0_outputs(3499) <= '1';
    layer0_outputs(3500) <= inputs(206);
    layer0_outputs(3501) <= (inputs(190)) and not (inputs(245));
    layer0_outputs(3502) <= not(inputs(4)) or (inputs(240));
    layer0_outputs(3503) <= inputs(83);
    layer0_outputs(3504) <= (inputs(205)) and (inputs(220));
    layer0_outputs(3505) <= not(inputs(8)) or (inputs(205));
    layer0_outputs(3506) <= inputs(32);
    layer0_outputs(3507) <= (inputs(104)) and not (inputs(51));
    layer0_outputs(3508) <= (inputs(56)) or (inputs(157));
    layer0_outputs(3509) <= (inputs(230)) and not (inputs(106));
    layer0_outputs(3510) <= (inputs(203)) or (inputs(141));
    layer0_outputs(3511) <= not((inputs(34)) or (inputs(199)));
    layer0_outputs(3512) <= not(inputs(173));
    layer0_outputs(3513) <= (inputs(183)) and not (inputs(53));
    layer0_outputs(3514) <= not((inputs(255)) or (inputs(85)));
    layer0_outputs(3515) <= not((inputs(33)) and (inputs(207)));
    layer0_outputs(3516) <= '1';
    layer0_outputs(3517) <= not(inputs(133)) or (inputs(211));
    layer0_outputs(3518) <= inputs(252);
    layer0_outputs(3519) <= not(inputs(248));
    layer0_outputs(3520) <= (inputs(76)) and not (inputs(128));
    layer0_outputs(3521) <= not(inputs(44)) or (inputs(223));
    layer0_outputs(3522) <= inputs(39);
    layer0_outputs(3523) <= not(inputs(61));
    layer0_outputs(3524) <= inputs(61);
    layer0_outputs(3525) <= inputs(99);
    layer0_outputs(3526) <= not((inputs(108)) and (inputs(84)));
    layer0_outputs(3527) <= (inputs(156)) or (inputs(172));
    layer0_outputs(3528) <= (inputs(208)) xor (inputs(35));
    layer0_outputs(3529) <= (inputs(60)) and not (inputs(120));
    layer0_outputs(3530) <= not((inputs(253)) xor (inputs(5)));
    layer0_outputs(3531) <= (inputs(48)) and not (inputs(55));
    layer0_outputs(3532) <= inputs(74);
    layer0_outputs(3533) <= not(inputs(20));
    layer0_outputs(3534) <= not(inputs(151));
    layer0_outputs(3535) <= (inputs(194)) and not (inputs(32));
    layer0_outputs(3536) <= (inputs(83)) and (inputs(92));
    layer0_outputs(3537) <= not(inputs(126));
    layer0_outputs(3538) <= (inputs(235)) and not (inputs(147));
    layer0_outputs(3539) <= not((inputs(64)) xor (inputs(84)));
    layer0_outputs(3540) <= inputs(182);
    layer0_outputs(3541) <= (inputs(157)) xor (inputs(126));
    layer0_outputs(3542) <= inputs(211);
    layer0_outputs(3543) <= (inputs(159)) xor (inputs(227));
    layer0_outputs(3544) <= not(inputs(41));
    layer0_outputs(3545) <= not(inputs(162)) or (inputs(130));
    layer0_outputs(3546) <= not(inputs(131));
    layer0_outputs(3547) <= not((inputs(98)) xor (inputs(177)));
    layer0_outputs(3548) <= not(inputs(248));
    layer0_outputs(3549) <= not(inputs(85));
    layer0_outputs(3550) <= (inputs(37)) and not (inputs(0));
    layer0_outputs(3551) <= not(inputs(151)) or (inputs(226));
    layer0_outputs(3552) <= not(inputs(25)) or (inputs(99));
    layer0_outputs(3553) <= '0';
    layer0_outputs(3554) <= (inputs(111)) xor (inputs(206));
    layer0_outputs(3555) <= (inputs(207)) and (inputs(47));
    layer0_outputs(3556) <= not((inputs(188)) xor (inputs(246)));
    layer0_outputs(3557) <= not(inputs(254));
    layer0_outputs(3558) <= not((inputs(24)) or (inputs(120)));
    layer0_outputs(3559) <= not(inputs(52)) or (inputs(156));
    layer0_outputs(3560) <= inputs(107);
    layer0_outputs(3561) <= (inputs(232)) and not (inputs(237));
    layer0_outputs(3562) <= '0';
    layer0_outputs(3563) <= inputs(104);
    layer0_outputs(3564) <= not(inputs(106));
    layer0_outputs(3565) <= (inputs(196)) or (inputs(126));
    layer0_outputs(3566) <= not(inputs(85)) or (inputs(139));
    layer0_outputs(3567) <= not(inputs(66));
    layer0_outputs(3568) <= (inputs(220)) and (inputs(250));
    layer0_outputs(3569) <= not((inputs(228)) or (inputs(160)));
    layer0_outputs(3570) <= (inputs(185)) and not (inputs(42));
    layer0_outputs(3571) <= (inputs(155)) or (inputs(35));
    layer0_outputs(3572) <= not(inputs(137)) or (inputs(188));
    layer0_outputs(3573) <= inputs(105);
    layer0_outputs(3574) <= inputs(234);
    layer0_outputs(3575) <= (inputs(88)) and not (inputs(211));
    layer0_outputs(3576) <= (inputs(154)) or (inputs(184));
    layer0_outputs(3577) <= inputs(107);
    layer0_outputs(3578) <= not(inputs(163)) or (inputs(235));
    layer0_outputs(3579) <= not((inputs(176)) and (inputs(50)));
    layer0_outputs(3580) <= not(inputs(206)) or (inputs(254));
    layer0_outputs(3581) <= not((inputs(20)) xor (inputs(78)));
    layer0_outputs(3582) <= (inputs(100)) and not (inputs(47));
    layer0_outputs(3583) <= not(inputs(225));
    layer0_outputs(3584) <= not(inputs(226));
    layer0_outputs(3585) <= inputs(114);
    layer0_outputs(3586) <= not(inputs(35));
    layer0_outputs(3587) <= not(inputs(117));
    layer0_outputs(3588) <= not(inputs(139)) or (inputs(112));
    layer0_outputs(3589) <= (inputs(230)) and (inputs(151));
    layer0_outputs(3590) <= (inputs(48)) and not (inputs(223));
    layer0_outputs(3591) <= not((inputs(112)) or (inputs(55)));
    layer0_outputs(3592) <= (inputs(10)) and not (inputs(127));
    layer0_outputs(3593) <= inputs(181);
    layer0_outputs(3594) <= inputs(169);
    layer0_outputs(3595) <= not(inputs(198));
    layer0_outputs(3596) <= not((inputs(232)) xor (inputs(184)));
    layer0_outputs(3597) <= not(inputs(91));
    layer0_outputs(3598) <= not(inputs(106));
    layer0_outputs(3599) <= (inputs(28)) and not (inputs(160));
    layer0_outputs(3600) <= (inputs(240)) or (inputs(166));
    layer0_outputs(3601) <= not((inputs(55)) xor (inputs(9)));
    layer0_outputs(3602) <= not((inputs(193)) xor (inputs(192)));
    layer0_outputs(3603) <= (inputs(127)) or (inputs(52));
    layer0_outputs(3604) <= (inputs(135)) and not (inputs(52));
    layer0_outputs(3605) <= (inputs(160)) or (inputs(162));
    layer0_outputs(3606) <= (inputs(252)) or (inputs(145));
    layer0_outputs(3607) <= not((inputs(123)) or (inputs(228)));
    layer0_outputs(3608) <= (inputs(224)) xor (inputs(247));
    layer0_outputs(3609) <= (inputs(126)) xor (inputs(156));
    layer0_outputs(3610) <= (inputs(73)) and (inputs(41));
    layer0_outputs(3611) <= inputs(200);
    layer0_outputs(3612) <= (inputs(132)) and not (inputs(83));
    layer0_outputs(3613) <= (inputs(107)) xor (inputs(156));
    layer0_outputs(3614) <= not(inputs(86));
    layer0_outputs(3615) <= '0';
    layer0_outputs(3616) <= not(inputs(251));
    layer0_outputs(3617) <= not((inputs(27)) or (inputs(204)));
    layer0_outputs(3618) <= '1';
    layer0_outputs(3619) <= not((inputs(178)) or (inputs(192)));
    layer0_outputs(3620) <= (inputs(193)) and not (inputs(253));
    layer0_outputs(3621) <= inputs(126);
    layer0_outputs(3622) <= inputs(29);
    layer0_outputs(3623) <= not((inputs(54)) and (inputs(194)));
    layer0_outputs(3624) <= inputs(1);
    layer0_outputs(3625) <= not(inputs(15)) or (inputs(17));
    layer0_outputs(3626) <= not((inputs(90)) xor (inputs(31)));
    layer0_outputs(3627) <= not(inputs(38));
    layer0_outputs(3628) <= not((inputs(91)) xor (inputs(124)));
    layer0_outputs(3629) <= (inputs(210)) or (inputs(194));
    layer0_outputs(3630) <= not(inputs(144));
    layer0_outputs(3631) <= not(inputs(130));
    layer0_outputs(3632) <= (inputs(107)) and not (inputs(172));
    layer0_outputs(3633) <= not(inputs(194));
    layer0_outputs(3634) <= inputs(200);
    layer0_outputs(3635) <= (inputs(183)) and not (inputs(201));
    layer0_outputs(3636) <= (inputs(252)) or (inputs(77));
    layer0_outputs(3637) <= not(inputs(0));
    layer0_outputs(3638) <= not((inputs(252)) or (inputs(182)));
    layer0_outputs(3639) <= (inputs(143)) and (inputs(55));
    layer0_outputs(3640) <= inputs(76);
    layer0_outputs(3641) <= not(inputs(3));
    layer0_outputs(3642) <= not(inputs(46)) or (inputs(123));
    layer0_outputs(3643) <= (inputs(42)) or (inputs(93));
    layer0_outputs(3644) <= inputs(82);
    layer0_outputs(3645) <= (inputs(83)) xor (inputs(117));
    layer0_outputs(3646) <= not(inputs(117));
    layer0_outputs(3647) <= inputs(232);
    layer0_outputs(3648) <= not(inputs(149));
    layer0_outputs(3649) <= not((inputs(161)) and (inputs(196)));
    layer0_outputs(3650) <= (inputs(147)) or (inputs(80));
    layer0_outputs(3651) <= not(inputs(235));
    layer0_outputs(3652) <= not(inputs(131));
    layer0_outputs(3653) <= (inputs(104)) and not (inputs(109));
    layer0_outputs(3654) <= (inputs(205)) xor (inputs(140));
    layer0_outputs(3655) <= not(inputs(41));
    layer0_outputs(3656) <= (inputs(205)) and (inputs(67));
    layer0_outputs(3657) <= inputs(236);
    layer0_outputs(3658) <= inputs(29);
    layer0_outputs(3659) <= (inputs(69)) or (inputs(28));
    layer0_outputs(3660) <= (inputs(243)) xor (inputs(142));
    layer0_outputs(3661) <= not(inputs(237)) or (inputs(125));
    layer0_outputs(3662) <= inputs(207);
    layer0_outputs(3663) <= (inputs(156)) or (inputs(196));
    layer0_outputs(3664) <= not(inputs(232));
    layer0_outputs(3665) <= (inputs(178)) or (inputs(117));
    layer0_outputs(3666) <= (inputs(88)) or (inputs(19));
    layer0_outputs(3667) <= (inputs(1)) or (inputs(235));
    layer0_outputs(3668) <= (inputs(208)) or (inputs(24));
    layer0_outputs(3669) <= (inputs(251)) and (inputs(199));
    layer0_outputs(3670) <= inputs(106);
    layer0_outputs(3671) <= (inputs(103)) and not (inputs(148));
    layer0_outputs(3672) <= not(inputs(116)) or (inputs(200));
    layer0_outputs(3673) <= (inputs(82)) and not (inputs(127));
    layer0_outputs(3674) <= not(inputs(49)) or (inputs(133));
    layer0_outputs(3675) <= (inputs(178)) and not (inputs(249));
    layer0_outputs(3676) <= (inputs(47)) xor (inputs(65));
    layer0_outputs(3677) <= '0';
    layer0_outputs(3678) <= (inputs(118)) and not (inputs(48));
    layer0_outputs(3679) <= not((inputs(201)) or (inputs(19)));
    layer0_outputs(3680) <= not((inputs(150)) or (inputs(122)));
    layer0_outputs(3681) <= (inputs(108)) xor (inputs(175));
    layer0_outputs(3682) <= not(inputs(181));
    layer0_outputs(3683) <= not((inputs(211)) or (inputs(129)));
    layer0_outputs(3684) <= not((inputs(7)) or (inputs(70)));
    layer0_outputs(3685) <= inputs(177);
    layer0_outputs(3686) <= (inputs(78)) or (inputs(26));
    layer0_outputs(3687) <= (inputs(55)) and (inputs(72));
    layer0_outputs(3688) <= (inputs(37)) and not (inputs(190));
    layer0_outputs(3689) <= not(inputs(210));
    layer0_outputs(3690) <= inputs(73);
    layer0_outputs(3691) <= '1';
    layer0_outputs(3692) <= not(inputs(93));
    layer0_outputs(3693) <= not(inputs(7)) or (inputs(145));
    layer0_outputs(3694) <= (inputs(29)) or (inputs(149));
    layer0_outputs(3695) <= '1';
    layer0_outputs(3696) <= not(inputs(113));
    layer0_outputs(3697) <= inputs(150);
    layer0_outputs(3698) <= (inputs(98)) and not (inputs(1));
    layer0_outputs(3699) <= not(inputs(156));
    layer0_outputs(3700) <= (inputs(68)) or (inputs(7));
    layer0_outputs(3701) <= (inputs(48)) xor (inputs(76));
    layer0_outputs(3702) <= (inputs(184)) or (inputs(183));
    layer0_outputs(3703) <= not(inputs(83)) or (inputs(153));
    layer0_outputs(3704) <= (inputs(224)) and not (inputs(143));
    layer0_outputs(3705) <= '1';
    layer0_outputs(3706) <= (inputs(215)) and (inputs(212));
    layer0_outputs(3707) <= (inputs(53)) and (inputs(37));
    layer0_outputs(3708) <= (inputs(235)) xor (inputs(171));
    layer0_outputs(3709) <= not(inputs(90));
    layer0_outputs(3710) <= (inputs(221)) or (inputs(147));
    layer0_outputs(3711) <= inputs(251);
    layer0_outputs(3712) <= not(inputs(25));
    layer0_outputs(3713) <= inputs(166);
    layer0_outputs(3714) <= '1';
    layer0_outputs(3715) <= (inputs(69)) or (inputs(112));
    layer0_outputs(3716) <= not((inputs(92)) xor (inputs(87)));
    layer0_outputs(3717) <= (inputs(222)) or (inputs(194));
    layer0_outputs(3718) <= (inputs(58)) and not (inputs(150));
    layer0_outputs(3719) <= not(inputs(28)) or (inputs(116));
    layer0_outputs(3720) <= (inputs(210)) or (inputs(117));
    layer0_outputs(3721) <= not(inputs(88)) or (inputs(80));
    layer0_outputs(3722) <= (inputs(168)) and not (inputs(95));
    layer0_outputs(3723) <= not(inputs(102)) or (inputs(67));
    layer0_outputs(3724) <= inputs(8);
    layer0_outputs(3725) <= not((inputs(89)) and (inputs(65)));
    layer0_outputs(3726) <= not(inputs(185));
    layer0_outputs(3727) <= not(inputs(186));
    layer0_outputs(3728) <= (inputs(232)) and not (inputs(130));
    layer0_outputs(3729) <= not((inputs(44)) and (inputs(25)));
    layer0_outputs(3730) <= inputs(18);
    layer0_outputs(3731) <= inputs(54);
    layer0_outputs(3732) <= not((inputs(86)) xor (inputs(232)));
    layer0_outputs(3733) <= '1';
    layer0_outputs(3734) <= not((inputs(177)) or (inputs(252)));
    layer0_outputs(3735) <= inputs(214);
    layer0_outputs(3736) <= inputs(105);
    layer0_outputs(3737) <= (inputs(151)) and not (inputs(5));
    layer0_outputs(3738) <= not((inputs(29)) and (inputs(229)));
    layer0_outputs(3739) <= inputs(240);
    layer0_outputs(3740) <= not(inputs(151));
    layer0_outputs(3741) <= (inputs(198)) and not (inputs(113));
    layer0_outputs(3742) <= '1';
    layer0_outputs(3743) <= not(inputs(167));
    layer0_outputs(3744) <= inputs(229);
    layer0_outputs(3745) <= not((inputs(95)) or (inputs(39)));
    layer0_outputs(3746) <= (inputs(137)) or (inputs(250));
    layer0_outputs(3747) <= (inputs(170)) or (inputs(122));
    layer0_outputs(3748) <= not((inputs(18)) or (inputs(41)));
    layer0_outputs(3749) <= inputs(172);
    layer0_outputs(3750) <= not(inputs(53)) or (inputs(204));
    layer0_outputs(3751) <= (inputs(117)) or (inputs(221));
    layer0_outputs(3752) <= inputs(45);
    layer0_outputs(3753) <= not(inputs(48)) or (inputs(213));
    layer0_outputs(3754) <= not((inputs(107)) xor (inputs(45)));
    layer0_outputs(3755) <= not(inputs(178)) or (inputs(115));
    layer0_outputs(3756) <= not(inputs(38));
    layer0_outputs(3757) <= not(inputs(11)) or (inputs(32));
    layer0_outputs(3758) <= not(inputs(26));
    layer0_outputs(3759) <= not(inputs(93)) or (inputs(185));
    layer0_outputs(3760) <= (inputs(225)) or (inputs(104));
    layer0_outputs(3761) <= inputs(11);
    layer0_outputs(3762) <= not((inputs(192)) or (inputs(196)));
    layer0_outputs(3763) <= not(inputs(57));
    layer0_outputs(3764) <= (inputs(136)) and not (inputs(191));
    layer0_outputs(3765) <= not(inputs(126));
    layer0_outputs(3766) <= (inputs(181)) and not (inputs(201));
    layer0_outputs(3767) <= not((inputs(240)) or (inputs(29)));
    layer0_outputs(3768) <= (inputs(106)) and not (inputs(3));
    layer0_outputs(3769) <= not((inputs(28)) and (inputs(40)));
    layer0_outputs(3770) <= not(inputs(120));
    layer0_outputs(3771) <= not(inputs(184));
    layer0_outputs(3772) <= (inputs(222)) or (inputs(50));
    layer0_outputs(3773) <= inputs(212);
    layer0_outputs(3774) <= not(inputs(10)) or (inputs(219));
    layer0_outputs(3775) <= not((inputs(81)) xor (inputs(143)));
    layer0_outputs(3776) <= (inputs(179)) and not (inputs(193));
    layer0_outputs(3777) <= (inputs(239)) or (inputs(68));
    layer0_outputs(3778) <= not((inputs(8)) xor (inputs(203)));
    layer0_outputs(3779) <= not((inputs(194)) or (inputs(87)));
    layer0_outputs(3780) <= (inputs(25)) and not (inputs(192));
    layer0_outputs(3781) <= not(inputs(158));
    layer0_outputs(3782) <= not(inputs(87));
    layer0_outputs(3783) <= (inputs(230)) or (inputs(216));
    layer0_outputs(3784) <= not((inputs(219)) or (inputs(239)));
    layer0_outputs(3785) <= inputs(77);
    layer0_outputs(3786) <= (inputs(121)) and not (inputs(239));
    layer0_outputs(3787) <= inputs(62);
    layer0_outputs(3788) <= not(inputs(67));
    layer0_outputs(3789) <= inputs(158);
    layer0_outputs(3790) <= (inputs(158)) or (inputs(96));
    layer0_outputs(3791) <= not((inputs(119)) or (inputs(227)));
    layer0_outputs(3792) <= (inputs(192)) or (inputs(193));
    layer0_outputs(3793) <= inputs(93);
    layer0_outputs(3794) <= '0';
    layer0_outputs(3795) <= not((inputs(243)) and (inputs(9)));
    layer0_outputs(3796) <= inputs(31);
    layer0_outputs(3797) <= inputs(37);
    layer0_outputs(3798) <= not(inputs(107));
    layer0_outputs(3799) <= inputs(132);
    layer0_outputs(3800) <= not((inputs(196)) or (inputs(181)));
    layer0_outputs(3801) <= (inputs(157)) xor (inputs(251));
    layer0_outputs(3802) <= not(inputs(81)) or (inputs(95));
    layer0_outputs(3803) <= not(inputs(132));
    layer0_outputs(3804) <= inputs(113);
    layer0_outputs(3805) <= not((inputs(174)) or (inputs(17)));
    layer0_outputs(3806) <= not((inputs(9)) or (inputs(209)));
    layer0_outputs(3807) <= (inputs(99)) or (inputs(153));
    layer0_outputs(3808) <= inputs(237);
    layer0_outputs(3809) <= inputs(91);
    layer0_outputs(3810) <= not(inputs(103)) or (inputs(80));
    layer0_outputs(3811) <= not(inputs(173)) or (inputs(146));
    layer0_outputs(3812) <= '0';
    layer0_outputs(3813) <= not(inputs(217));
    layer0_outputs(3814) <= not(inputs(166));
    layer0_outputs(3815) <= (inputs(54)) and not (inputs(111));
    layer0_outputs(3816) <= not(inputs(176));
    layer0_outputs(3817) <= not(inputs(137)) or (inputs(97));
    layer0_outputs(3818) <= (inputs(127)) and not (inputs(255));
    layer0_outputs(3819) <= not((inputs(145)) or (inputs(187)));
    layer0_outputs(3820) <= inputs(135);
    layer0_outputs(3821) <= '0';
    layer0_outputs(3822) <= not((inputs(181)) or (inputs(65)));
    layer0_outputs(3823) <= not(inputs(60));
    layer0_outputs(3824) <= not((inputs(13)) xor (inputs(144)));
    layer0_outputs(3825) <= (inputs(79)) or (inputs(97));
    layer0_outputs(3826) <= (inputs(167)) and not (inputs(114));
    layer0_outputs(3827) <= (inputs(34)) and not (inputs(112));
    layer0_outputs(3828) <= (inputs(132)) and not (inputs(14));
    layer0_outputs(3829) <= '1';
    layer0_outputs(3830) <= '1';
    layer0_outputs(3831) <= not(inputs(221));
    layer0_outputs(3832) <= not((inputs(231)) or (inputs(115)));
    layer0_outputs(3833) <= (inputs(135)) and not (inputs(125));
    layer0_outputs(3834) <= inputs(90);
    layer0_outputs(3835) <= not(inputs(195));
    layer0_outputs(3836) <= not(inputs(25)) or (inputs(229));
    layer0_outputs(3837) <= '1';
    layer0_outputs(3838) <= '0';
    layer0_outputs(3839) <= not((inputs(81)) xor (inputs(176)));
    layer0_outputs(3840) <= '0';
    layer0_outputs(3841) <= not((inputs(59)) or (inputs(51)));
    layer0_outputs(3842) <= not((inputs(102)) or (inputs(87)));
    layer0_outputs(3843) <= (inputs(58)) and (inputs(81));
    layer0_outputs(3844) <= (inputs(87)) xor (inputs(43));
    layer0_outputs(3845) <= (inputs(123)) xor (inputs(175));
    layer0_outputs(3846) <= '1';
    layer0_outputs(3847) <= (inputs(173)) and not (inputs(137));
    layer0_outputs(3848) <= not((inputs(13)) xor (inputs(225)));
    layer0_outputs(3849) <= inputs(104);
    layer0_outputs(3850) <= not(inputs(142)) or (inputs(153));
    layer0_outputs(3851) <= (inputs(185)) and (inputs(246));
    layer0_outputs(3852) <= not(inputs(188));
    layer0_outputs(3853) <= not(inputs(119));
    layer0_outputs(3854) <= (inputs(49)) and not (inputs(203));
    layer0_outputs(3855) <= inputs(134);
    layer0_outputs(3856) <= inputs(8);
    layer0_outputs(3857) <= (inputs(131)) or (inputs(145));
    layer0_outputs(3858) <= (inputs(109)) or (inputs(215));
    layer0_outputs(3859) <= not((inputs(70)) and (inputs(225)));
    layer0_outputs(3860) <= not(inputs(140));
    layer0_outputs(3861) <= '0';
    layer0_outputs(3862) <= (inputs(165)) or (inputs(209));
    layer0_outputs(3863) <= (inputs(113)) xor (inputs(219));
    layer0_outputs(3864) <= inputs(107);
    layer0_outputs(3865) <= (inputs(184)) and not (inputs(142));
    layer0_outputs(3866) <= not((inputs(199)) and (inputs(182)));
    layer0_outputs(3867) <= inputs(229);
    layer0_outputs(3868) <= (inputs(0)) and not (inputs(183));
    layer0_outputs(3869) <= not(inputs(29));
    layer0_outputs(3870) <= not((inputs(195)) xor (inputs(33)));
    layer0_outputs(3871) <= '1';
    layer0_outputs(3872) <= not(inputs(91));
    layer0_outputs(3873) <= not(inputs(162)) or (inputs(54));
    layer0_outputs(3874) <= not(inputs(246)) or (inputs(148));
    layer0_outputs(3875) <= (inputs(78)) or (inputs(101));
    layer0_outputs(3876) <= (inputs(72)) or (inputs(14));
    layer0_outputs(3877) <= not((inputs(68)) and (inputs(27)));
    layer0_outputs(3878) <= inputs(207);
    layer0_outputs(3879) <= not((inputs(175)) or (inputs(86)));
    layer0_outputs(3880) <= inputs(41);
    layer0_outputs(3881) <= (inputs(195)) and not (inputs(91));
    layer0_outputs(3882) <= (inputs(151)) and not (inputs(91));
    layer0_outputs(3883) <= inputs(123);
    layer0_outputs(3884) <= (inputs(139)) and not (inputs(68));
    layer0_outputs(3885) <= (inputs(159)) and not (inputs(207));
    layer0_outputs(3886) <= not(inputs(154)) or (inputs(191));
    layer0_outputs(3887) <= inputs(157);
    layer0_outputs(3888) <= inputs(105);
    layer0_outputs(3889) <= '0';
    layer0_outputs(3890) <= inputs(202);
    layer0_outputs(3891) <= (inputs(162)) xor (inputs(133));
    layer0_outputs(3892) <= '0';
    layer0_outputs(3893) <= (inputs(33)) or (inputs(91));
    layer0_outputs(3894) <= (inputs(243)) and not (inputs(52));
    layer0_outputs(3895) <= not(inputs(163));
    layer0_outputs(3896) <= inputs(134);
    layer0_outputs(3897) <= (inputs(30)) and (inputs(231));
    layer0_outputs(3898) <= (inputs(172)) and not (inputs(14));
    layer0_outputs(3899) <= not((inputs(119)) or (inputs(223)));
    layer0_outputs(3900) <= (inputs(183)) and not (inputs(248));
    layer0_outputs(3901) <= not(inputs(25)) or (inputs(86));
    layer0_outputs(3902) <= inputs(131);
    layer0_outputs(3903) <= (inputs(117)) or (inputs(194));
    layer0_outputs(3904) <= not((inputs(50)) or (inputs(60)));
    layer0_outputs(3905) <= not((inputs(12)) xor (inputs(33)));
    layer0_outputs(3906) <= (inputs(62)) or (inputs(106));
    layer0_outputs(3907) <= not(inputs(143));
    layer0_outputs(3908) <= not(inputs(61)) or (inputs(229));
    layer0_outputs(3909) <= not(inputs(177));
    layer0_outputs(3910) <= not(inputs(234));
    layer0_outputs(3911) <= not((inputs(63)) or (inputs(38)));
    layer0_outputs(3912) <= not(inputs(46));
    layer0_outputs(3913) <= inputs(89);
    layer0_outputs(3914) <= not(inputs(94));
    layer0_outputs(3915) <= not(inputs(90)) or (inputs(220));
    layer0_outputs(3916) <= (inputs(142)) or (inputs(248));
    layer0_outputs(3917) <= not(inputs(219)) or (inputs(31));
    layer0_outputs(3918) <= inputs(71);
    layer0_outputs(3919) <= '1';
    layer0_outputs(3920) <= (inputs(112)) and not (inputs(236));
    layer0_outputs(3921) <= inputs(123);
    layer0_outputs(3922) <= not((inputs(140)) or (inputs(1)));
    layer0_outputs(3923) <= inputs(2);
    layer0_outputs(3924) <= (inputs(160)) or (inputs(62));
    layer0_outputs(3925) <= not(inputs(239)) or (inputs(134));
    layer0_outputs(3926) <= not(inputs(24)) or (inputs(219));
    layer0_outputs(3927) <= inputs(77);
    layer0_outputs(3928) <= inputs(120);
    layer0_outputs(3929) <= not(inputs(221)) or (inputs(125));
    layer0_outputs(3930) <= (inputs(233)) and not (inputs(20));
    layer0_outputs(3931) <= not(inputs(156));
    layer0_outputs(3932) <= inputs(175);
    layer0_outputs(3933) <= not(inputs(127)) or (inputs(224));
    layer0_outputs(3934) <= '1';
    layer0_outputs(3935) <= (inputs(121)) or (inputs(41));
    layer0_outputs(3936) <= (inputs(182)) and (inputs(90));
    layer0_outputs(3937) <= not(inputs(79)) or (inputs(31));
    layer0_outputs(3938) <= (inputs(2)) and not (inputs(76));
    layer0_outputs(3939) <= (inputs(133)) and not (inputs(1));
    layer0_outputs(3940) <= not(inputs(110)) or (inputs(16));
    layer0_outputs(3941) <= not((inputs(184)) xor (inputs(255)));
    layer0_outputs(3942) <= not((inputs(125)) or (inputs(100)));
    layer0_outputs(3943) <= not((inputs(18)) or (inputs(17)));
    layer0_outputs(3944) <= (inputs(216)) and not (inputs(31));
    layer0_outputs(3945) <= inputs(118);
    layer0_outputs(3946) <= not((inputs(66)) and (inputs(26)));
    layer0_outputs(3947) <= inputs(47);
    layer0_outputs(3948) <= (inputs(172)) and not (inputs(222));
    layer0_outputs(3949) <= not(inputs(10)) or (inputs(160));
    layer0_outputs(3950) <= (inputs(21)) and not (inputs(94));
    layer0_outputs(3951) <= inputs(54);
    layer0_outputs(3952) <= (inputs(158)) and not (inputs(123));
    layer0_outputs(3953) <= not(inputs(231));
    layer0_outputs(3954) <= inputs(81);
    layer0_outputs(3955) <= not(inputs(26)) or (inputs(203));
    layer0_outputs(3956) <= inputs(109);
    layer0_outputs(3957) <= not((inputs(235)) or (inputs(19)));
    layer0_outputs(3958) <= not(inputs(22));
    layer0_outputs(3959) <= not(inputs(109));
    layer0_outputs(3960) <= inputs(25);
    layer0_outputs(3961) <= (inputs(109)) xor (inputs(181));
    layer0_outputs(3962) <= inputs(106);
    layer0_outputs(3963) <= not(inputs(25));
    layer0_outputs(3964) <= '1';
    layer0_outputs(3965) <= not(inputs(128));
    layer0_outputs(3966) <= inputs(74);
    layer0_outputs(3967) <= (inputs(75)) and not (inputs(242));
    layer0_outputs(3968) <= not((inputs(47)) or (inputs(22)));
    layer0_outputs(3969) <= inputs(14);
    layer0_outputs(3970) <= (inputs(129)) or (inputs(213));
    layer0_outputs(3971) <= (inputs(58)) or (inputs(66));
    layer0_outputs(3972) <= not(inputs(61));
    layer0_outputs(3973) <= inputs(40);
    layer0_outputs(3974) <= not((inputs(87)) or (inputs(218)));
    layer0_outputs(3975) <= inputs(225);
    layer0_outputs(3976) <= (inputs(78)) xor (inputs(4));
    layer0_outputs(3977) <= not(inputs(232)) or (inputs(103));
    layer0_outputs(3978) <= inputs(187);
    layer0_outputs(3979) <= (inputs(170)) and (inputs(74));
    layer0_outputs(3980) <= not((inputs(102)) or (inputs(50)));
    layer0_outputs(3981) <= inputs(178);
    layer0_outputs(3982) <= not((inputs(88)) or (inputs(160)));
    layer0_outputs(3983) <= (inputs(208)) and not (inputs(212));
    layer0_outputs(3984) <= not((inputs(138)) xor (inputs(217)));
    layer0_outputs(3985) <= not(inputs(182));
    layer0_outputs(3986) <= (inputs(60)) and not (inputs(152));
    layer0_outputs(3987) <= not(inputs(67)) or (inputs(179));
    layer0_outputs(3988) <= not((inputs(20)) and (inputs(34)));
    layer0_outputs(3989) <= (inputs(20)) xor (inputs(102));
    layer0_outputs(3990) <= inputs(150);
    layer0_outputs(3991) <= not((inputs(250)) or (inputs(81)));
    layer0_outputs(3992) <= (inputs(214)) and not (inputs(209));
    layer0_outputs(3993) <= (inputs(206)) and (inputs(124));
    layer0_outputs(3994) <= not((inputs(108)) or (inputs(83)));
    layer0_outputs(3995) <= inputs(51);
    layer0_outputs(3996) <= (inputs(43)) or (inputs(77));
    layer0_outputs(3997) <= not(inputs(229));
    layer0_outputs(3998) <= not(inputs(23)) or (inputs(201));
    layer0_outputs(3999) <= inputs(50);
    layer0_outputs(4000) <= not(inputs(173));
    layer0_outputs(4001) <= not((inputs(186)) xor (inputs(217)));
    layer0_outputs(4002) <= inputs(105);
    layer0_outputs(4003) <= '1';
    layer0_outputs(4004) <= not((inputs(4)) or (inputs(136)));
    layer0_outputs(4005) <= not((inputs(98)) xor (inputs(66)));
    layer0_outputs(4006) <= inputs(228);
    layer0_outputs(4007) <= not((inputs(108)) and (inputs(30)));
    layer0_outputs(4008) <= (inputs(44)) and not (inputs(140));
    layer0_outputs(4009) <= (inputs(180)) and not (inputs(88));
    layer0_outputs(4010) <= inputs(186);
    layer0_outputs(4011) <= '0';
    layer0_outputs(4012) <= not(inputs(19));
    layer0_outputs(4013) <= (inputs(47)) and not (inputs(64));
    layer0_outputs(4014) <= not(inputs(177)) or (inputs(189));
    layer0_outputs(4015) <= not(inputs(124));
    layer0_outputs(4016) <= not(inputs(70));
    layer0_outputs(4017) <= (inputs(58)) and not (inputs(173));
    layer0_outputs(4018) <= not((inputs(238)) xor (inputs(187)));
    layer0_outputs(4019) <= inputs(86);
    layer0_outputs(4020) <= '1';
    layer0_outputs(4021) <= (inputs(157)) and not (inputs(0));
    layer0_outputs(4022) <= (inputs(173)) or (inputs(93));
    layer0_outputs(4023) <= not(inputs(161));
    layer0_outputs(4024) <= not(inputs(38)) or (inputs(220));
    layer0_outputs(4025) <= (inputs(108)) or (inputs(99));
    layer0_outputs(4026) <= not(inputs(204)) or (inputs(97));
    layer0_outputs(4027) <= (inputs(4)) or (inputs(212));
    layer0_outputs(4028) <= not((inputs(224)) and (inputs(218)));
    layer0_outputs(4029) <= not(inputs(89));
    layer0_outputs(4030) <= (inputs(26)) or (inputs(45));
    layer0_outputs(4031) <= (inputs(46)) xor (inputs(218));
    layer0_outputs(4032) <= not((inputs(128)) or (inputs(145)));
    layer0_outputs(4033) <= not(inputs(100));
    layer0_outputs(4034) <= '0';
    layer0_outputs(4035) <= not((inputs(20)) or (inputs(206)));
    layer0_outputs(4036) <= (inputs(219)) and (inputs(120));
    layer0_outputs(4037) <= not(inputs(77)) or (inputs(102));
    layer0_outputs(4038) <= (inputs(121)) or (inputs(135));
    layer0_outputs(4039) <= inputs(94);
    layer0_outputs(4040) <= (inputs(57)) and not (inputs(112));
    layer0_outputs(4041) <= '0';
    layer0_outputs(4042) <= (inputs(152)) and not (inputs(73));
    layer0_outputs(4043) <= (inputs(32)) or (inputs(164));
    layer0_outputs(4044) <= (inputs(6)) and not (inputs(140));
    layer0_outputs(4045) <= not((inputs(115)) and (inputs(139)));
    layer0_outputs(4046) <= (inputs(87)) and not (inputs(66));
    layer0_outputs(4047) <= (inputs(186)) and not (inputs(33));
    layer0_outputs(4048) <= (inputs(167)) and not (inputs(79));
    layer0_outputs(4049) <= (inputs(201)) and not (inputs(18));
    layer0_outputs(4050) <= inputs(75);
    layer0_outputs(4051) <= not((inputs(75)) xor (inputs(195)));
    layer0_outputs(4052) <= not(inputs(90));
    layer0_outputs(4053) <= (inputs(61)) xor (inputs(30));
    layer0_outputs(4054) <= not(inputs(109)) or (inputs(130));
    layer0_outputs(4055) <= inputs(164);
    layer0_outputs(4056) <= (inputs(143)) and not (inputs(163));
    layer0_outputs(4057) <= (inputs(114)) or (inputs(84));
    layer0_outputs(4058) <= not(inputs(114));
    layer0_outputs(4059) <= not((inputs(244)) or (inputs(249)));
    layer0_outputs(4060) <= (inputs(55)) and not (inputs(103));
    layer0_outputs(4061) <= '0';
    layer0_outputs(4062) <= inputs(117);
    layer0_outputs(4063) <= inputs(22);
    layer0_outputs(4064) <= inputs(54);
    layer0_outputs(4065) <= not((inputs(158)) or (inputs(164)));
    layer0_outputs(4066) <= inputs(252);
    layer0_outputs(4067) <= (inputs(102)) and not (inputs(7));
    layer0_outputs(4068) <= '1';
    layer0_outputs(4069) <= inputs(82);
    layer0_outputs(4070) <= not(inputs(104)) or (inputs(143));
    layer0_outputs(4071) <= not(inputs(248));
    layer0_outputs(4072) <= (inputs(61)) and not (inputs(126));
    layer0_outputs(4073) <= (inputs(95)) and not (inputs(55));
    layer0_outputs(4074) <= inputs(85);
    layer0_outputs(4075) <= not((inputs(57)) and (inputs(21)));
    layer0_outputs(4076) <= (inputs(87)) and not (inputs(79));
    layer0_outputs(4077) <= not(inputs(187));
    layer0_outputs(4078) <= (inputs(199)) and not (inputs(155));
    layer0_outputs(4079) <= not(inputs(161));
    layer0_outputs(4080) <= (inputs(48)) and not (inputs(79));
    layer0_outputs(4081) <= (inputs(8)) xor (inputs(34));
    layer0_outputs(4082) <= (inputs(89)) and (inputs(21));
    layer0_outputs(4083) <= not(inputs(234)) or (inputs(241));
    layer0_outputs(4084) <= (inputs(86)) or (inputs(112));
    layer0_outputs(4085) <= (inputs(85)) and (inputs(29));
    layer0_outputs(4086) <= (inputs(117)) or (inputs(234));
    layer0_outputs(4087) <= not(inputs(245));
    layer0_outputs(4088) <= (inputs(66)) and (inputs(140));
    layer0_outputs(4089) <= (inputs(42)) and not (inputs(173));
    layer0_outputs(4090) <= (inputs(194)) or (inputs(234));
    layer0_outputs(4091) <= not(inputs(92));
    layer0_outputs(4092) <= not(inputs(37));
    layer0_outputs(4093) <= not(inputs(172)) or (inputs(9));
    layer0_outputs(4094) <= (inputs(244)) xor (inputs(173));
    layer0_outputs(4095) <= not((inputs(106)) xor (inputs(101)));
    layer0_outputs(4096) <= inputs(78);
    layer0_outputs(4097) <= (inputs(235)) or (inputs(85));
    layer0_outputs(4098) <= not(inputs(111)) or (inputs(48));
    layer0_outputs(4099) <= inputs(62);
    layer0_outputs(4100) <= (inputs(111)) or (inputs(248));
    layer0_outputs(4101) <= not(inputs(146));
    layer0_outputs(4102) <= (inputs(167)) or (inputs(64));
    layer0_outputs(4103) <= (inputs(230)) and not (inputs(108));
    layer0_outputs(4104) <= not(inputs(24));
    layer0_outputs(4105) <= (inputs(192)) and not (inputs(79));
    layer0_outputs(4106) <= (inputs(84)) and not (inputs(197));
    layer0_outputs(4107) <= inputs(104);
    layer0_outputs(4108) <= not((inputs(93)) or (inputs(254)));
    layer0_outputs(4109) <= not((inputs(99)) or (inputs(117)));
    layer0_outputs(4110) <= (inputs(18)) or (inputs(127));
    layer0_outputs(4111) <= not(inputs(35)) or (inputs(117));
    layer0_outputs(4112) <= (inputs(22)) xor (inputs(254));
    layer0_outputs(4113) <= (inputs(107)) or (inputs(62));
    layer0_outputs(4114) <= inputs(212);
    layer0_outputs(4115) <= inputs(230);
    layer0_outputs(4116) <= (inputs(24)) xor (inputs(48));
    layer0_outputs(4117) <= (inputs(237)) or (inputs(25));
    layer0_outputs(4118) <= not(inputs(182));
    layer0_outputs(4119) <= not(inputs(197));
    layer0_outputs(4120) <= not(inputs(252));
    layer0_outputs(4121) <= (inputs(222)) or (inputs(168));
    layer0_outputs(4122) <= not(inputs(112));
    layer0_outputs(4123) <= inputs(97);
    layer0_outputs(4124) <= (inputs(75)) and not (inputs(66));
    layer0_outputs(4125) <= (inputs(26)) xor (inputs(77));
    layer0_outputs(4126) <= not(inputs(117));
    layer0_outputs(4127) <= (inputs(230)) and (inputs(167));
    layer0_outputs(4128) <= (inputs(216)) and (inputs(51));
    layer0_outputs(4129) <= inputs(44);
    layer0_outputs(4130) <= not(inputs(108)) or (inputs(220));
    layer0_outputs(4131) <= inputs(224);
    layer0_outputs(4132) <= (inputs(226)) and not (inputs(254));
    layer0_outputs(4133) <= not(inputs(100)) or (inputs(165));
    layer0_outputs(4134) <= not((inputs(109)) xor (inputs(219)));
    layer0_outputs(4135) <= (inputs(152)) and (inputs(11));
    layer0_outputs(4136) <= (inputs(171)) and not (inputs(12));
    layer0_outputs(4137) <= inputs(136);
    layer0_outputs(4138) <= (inputs(39)) or (inputs(62));
    layer0_outputs(4139) <= inputs(190);
    layer0_outputs(4140) <= not(inputs(143)) or (inputs(158));
    layer0_outputs(4141) <= not(inputs(78)) or (inputs(46));
    layer0_outputs(4142) <= (inputs(172)) or (inputs(143));
    layer0_outputs(4143) <= not((inputs(174)) xor (inputs(86)));
    layer0_outputs(4144) <= not((inputs(159)) or (inputs(141)));
    layer0_outputs(4145) <= not((inputs(198)) xor (inputs(81)));
    layer0_outputs(4146) <= inputs(153);
    layer0_outputs(4147) <= inputs(89);
    layer0_outputs(4148) <= (inputs(189)) and not (inputs(37));
    layer0_outputs(4149) <= not(inputs(69));
    layer0_outputs(4150) <= not((inputs(184)) or (inputs(125)));
    layer0_outputs(4151) <= inputs(100);
    layer0_outputs(4152) <= not(inputs(63));
    layer0_outputs(4153) <= not(inputs(37));
    layer0_outputs(4154) <= (inputs(95)) xor (inputs(108));
    layer0_outputs(4155) <= inputs(8);
    layer0_outputs(4156) <= inputs(85);
    layer0_outputs(4157) <= inputs(93);
    layer0_outputs(4158) <= not(inputs(201));
    layer0_outputs(4159) <= not(inputs(161));
    layer0_outputs(4160) <= not((inputs(28)) or (inputs(115)));
    layer0_outputs(4161) <= not((inputs(112)) xor (inputs(48)));
    layer0_outputs(4162) <= (inputs(136)) and not (inputs(142));
    layer0_outputs(4163) <= (inputs(163)) and not (inputs(124));
    layer0_outputs(4164) <= not(inputs(150)) or (inputs(244));
    layer0_outputs(4165) <= not((inputs(113)) or (inputs(29)));
    layer0_outputs(4166) <= (inputs(175)) xor (inputs(222));
    layer0_outputs(4167) <= not(inputs(164));
    layer0_outputs(4168) <= not((inputs(164)) or (inputs(1)));
    layer0_outputs(4169) <= not(inputs(121));
    layer0_outputs(4170) <= (inputs(66)) and not (inputs(245));
    layer0_outputs(4171) <= not(inputs(233));
    layer0_outputs(4172) <= (inputs(7)) xor (inputs(224));
    layer0_outputs(4173) <= (inputs(205)) and not (inputs(206));
    layer0_outputs(4174) <= inputs(208);
    layer0_outputs(4175) <= not((inputs(5)) or (inputs(46)));
    layer0_outputs(4176) <= (inputs(95)) or (inputs(113));
    layer0_outputs(4177) <= inputs(174);
    layer0_outputs(4178) <= inputs(9);
    layer0_outputs(4179) <= inputs(111);
    layer0_outputs(4180) <= inputs(196);
    layer0_outputs(4181) <= inputs(60);
    layer0_outputs(4182) <= (inputs(21)) and not (inputs(199));
    layer0_outputs(4183) <= (inputs(21)) xor (inputs(67));
    layer0_outputs(4184) <= (inputs(69)) xor (inputs(98));
    layer0_outputs(4185) <= not(inputs(118)) or (inputs(235));
    layer0_outputs(4186) <= (inputs(184)) or (inputs(83));
    layer0_outputs(4187) <= (inputs(85)) xor (inputs(70));
    layer0_outputs(4188) <= (inputs(62)) xor (inputs(117));
    layer0_outputs(4189) <= not(inputs(70));
    layer0_outputs(4190) <= inputs(165);
    layer0_outputs(4191) <= not(inputs(210));
    layer0_outputs(4192) <= not(inputs(130)) or (inputs(161));
    layer0_outputs(4193) <= not(inputs(133)) or (inputs(158));
    layer0_outputs(4194) <= inputs(68);
    layer0_outputs(4195) <= (inputs(175)) and not (inputs(153));
    layer0_outputs(4196) <= '1';
    layer0_outputs(4197) <= inputs(89);
    layer0_outputs(4198) <= not((inputs(170)) xor (inputs(23)));
    layer0_outputs(4199) <= not(inputs(22));
    layer0_outputs(4200) <= (inputs(68)) xor (inputs(140));
    layer0_outputs(4201) <= inputs(138);
    layer0_outputs(4202) <= inputs(249);
    layer0_outputs(4203) <= not(inputs(236));
    layer0_outputs(4204) <= not((inputs(56)) or (inputs(72)));
    layer0_outputs(4205) <= inputs(12);
    layer0_outputs(4206) <= not(inputs(71));
    layer0_outputs(4207) <= inputs(163);
    layer0_outputs(4208) <= not((inputs(68)) or (inputs(109)));
    layer0_outputs(4209) <= (inputs(83)) and not (inputs(254));
    layer0_outputs(4210) <= inputs(93);
    layer0_outputs(4211) <= (inputs(173)) or (inputs(114));
    layer0_outputs(4212) <= not(inputs(155)) or (inputs(235));
    layer0_outputs(4213) <= not(inputs(101));
    layer0_outputs(4214) <= inputs(214);
    layer0_outputs(4215) <= not(inputs(211));
    layer0_outputs(4216) <= inputs(245);
    layer0_outputs(4217) <= not(inputs(187)) or (inputs(96));
    layer0_outputs(4218) <= (inputs(132)) xor (inputs(9));
    layer0_outputs(4219) <= inputs(163);
    layer0_outputs(4220) <= not(inputs(75));
    layer0_outputs(4221) <= not(inputs(167));
    layer0_outputs(4222) <= not((inputs(202)) and (inputs(189)));
    layer0_outputs(4223) <= not(inputs(152));
    layer0_outputs(4224) <= '1';
    layer0_outputs(4225) <= not(inputs(230));
    layer0_outputs(4226) <= inputs(35);
    layer0_outputs(4227) <= not((inputs(136)) xor (inputs(167)));
    layer0_outputs(4228) <= not(inputs(111)) or (inputs(237));
    layer0_outputs(4229) <= not((inputs(207)) xor (inputs(199)));
    layer0_outputs(4230) <= not(inputs(32)) or (inputs(229));
    layer0_outputs(4231) <= not(inputs(248)) or (inputs(77));
    layer0_outputs(4232) <= (inputs(126)) and not (inputs(40));
    layer0_outputs(4233) <= (inputs(131)) or (inputs(247));
    layer0_outputs(4234) <= not(inputs(159));
    layer0_outputs(4235) <= (inputs(64)) or (inputs(73));
    layer0_outputs(4236) <= not(inputs(166)) or (inputs(160));
    layer0_outputs(4237) <= (inputs(57)) or (inputs(179));
    layer0_outputs(4238) <= not(inputs(138));
    layer0_outputs(4239) <= inputs(19);
    layer0_outputs(4240) <= not(inputs(7));
    layer0_outputs(4241) <= (inputs(172)) or (inputs(28));
    layer0_outputs(4242) <= not(inputs(239));
    layer0_outputs(4243) <= not(inputs(17)) or (inputs(112));
    layer0_outputs(4244) <= (inputs(238)) xor (inputs(177));
    layer0_outputs(4245) <= inputs(54);
    layer0_outputs(4246) <= not(inputs(221));
    layer0_outputs(4247) <= inputs(220);
    layer0_outputs(4248) <= inputs(66);
    layer0_outputs(4249) <= '0';
    layer0_outputs(4250) <= (inputs(188)) xor (inputs(122));
    layer0_outputs(4251) <= '0';
    layer0_outputs(4252) <= not((inputs(150)) or (inputs(191)));
    layer0_outputs(4253) <= (inputs(115)) xor (inputs(103));
    layer0_outputs(4254) <= inputs(169);
    layer0_outputs(4255) <= not(inputs(56)) or (inputs(219));
    layer0_outputs(4256) <= inputs(77);
    layer0_outputs(4257) <= not((inputs(33)) or (inputs(121)));
    layer0_outputs(4258) <= not(inputs(148)) or (inputs(192));
    layer0_outputs(4259) <= inputs(246);
    layer0_outputs(4260) <= not((inputs(199)) xor (inputs(244)));
    layer0_outputs(4261) <= not(inputs(11));
    layer0_outputs(4262) <= (inputs(66)) xor (inputs(217));
    layer0_outputs(4263) <= (inputs(102)) and (inputs(183));
    layer0_outputs(4264) <= '0';
    layer0_outputs(4265) <= not(inputs(145));
    layer0_outputs(4266) <= (inputs(239)) and not (inputs(252));
    layer0_outputs(4267) <= not(inputs(192)) or (inputs(248));
    layer0_outputs(4268) <= not(inputs(172));
    layer0_outputs(4269) <= not(inputs(236));
    layer0_outputs(4270) <= inputs(100);
    layer0_outputs(4271) <= '0';
    layer0_outputs(4272) <= inputs(83);
    layer0_outputs(4273) <= (inputs(110)) xor (inputs(220));
    layer0_outputs(4274) <= not((inputs(204)) or (inputs(130)));
    layer0_outputs(4275) <= '1';
    layer0_outputs(4276) <= not(inputs(95));
    layer0_outputs(4277) <= not(inputs(78)) or (inputs(35));
    layer0_outputs(4278) <= not(inputs(58));
    layer0_outputs(4279) <= (inputs(226)) xor (inputs(16));
    layer0_outputs(4280) <= not((inputs(25)) xor (inputs(50)));
    layer0_outputs(4281) <= not(inputs(39));
    layer0_outputs(4282) <= not(inputs(44));
    layer0_outputs(4283) <= inputs(167);
    layer0_outputs(4284) <= (inputs(243)) and not (inputs(37));
    layer0_outputs(4285) <= (inputs(65)) and not (inputs(59));
    layer0_outputs(4286) <= (inputs(59)) or (inputs(120));
    layer0_outputs(4287) <= inputs(61);
    layer0_outputs(4288) <= (inputs(202)) or (inputs(111));
    layer0_outputs(4289) <= not((inputs(99)) or (inputs(243)));
    layer0_outputs(4290) <= (inputs(246)) or (inputs(21));
    layer0_outputs(4291) <= not((inputs(111)) or (inputs(75)));
    layer0_outputs(4292) <= (inputs(173)) or (inputs(53));
    layer0_outputs(4293) <= inputs(206);
    layer0_outputs(4294) <= not((inputs(140)) or (inputs(90)));
    layer0_outputs(4295) <= not((inputs(74)) or (inputs(35)));
    layer0_outputs(4296) <= not((inputs(14)) or (inputs(132)));
    layer0_outputs(4297) <= not(inputs(206));
    layer0_outputs(4298) <= (inputs(249)) and not (inputs(200));
    layer0_outputs(4299) <= not(inputs(20));
    layer0_outputs(4300) <= not(inputs(249)) or (inputs(143));
    layer0_outputs(4301) <= (inputs(196)) and not (inputs(203));
    layer0_outputs(4302) <= '0';
    layer0_outputs(4303) <= not(inputs(201));
    layer0_outputs(4304) <= (inputs(184)) or (inputs(243));
    layer0_outputs(4305) <= inputs(35);
    layer0_outputs(4306) <= inputs(29);
    layer0_outputs(4307) <= (inputs(61)) or (inputs(227));
    layer0_outputs(4308) <= not(inputs(237)) or (inputs(49));
    layer0_outputs(4309) <= inputs(5);
    layer0_outputs(4310) <= not((inputs(19)) or (inputs(37)));
    layer0_outputs(4311) <= (inputs(222)) xor (inputs(228));
    layer0_outputs(4312) <= not(inputs(29));
    layer0_outputs(4313) <= inputs(67);
    layer0_outputs(4314) <= '0';
    layer0_outputs(4315) <= not(inputs(134));
    layer0_outputs(4316) <= not((inputs(33)) and (inputs(12)));
    layer0_outputs(4317) <= not((inputs(60)) or (inputs(5)));
    layer0_outputs(4318) <= not((inputs(171)) or (inputs(144)));
    layer0_outputs(4319) <= not(inputs(117)) or (inputs(255));
    layer0_outputs(4320) <= not(inputs(122)) or (inputs(102));
    layer0_outputs(4321) <= not(inputs(248));
    layer0_outputs(4322) <= (inputs(93)) xor (inputs(183));
    layer0_outputs(4323) <= not(inputs(190));
    layer0_outputs(4324) <= inputs(42);
    layer0_outputs(4325) <= not((inputs(82)) or (inputs(196)));
    layer0_outputs(4326) <= not(inputs(242));
    layer0_outputs(4327) <= not(inputs(189)) or (inputs(31));
    layer0_outputs(4328) <= (inputs(34)) or (inputs(103));
    layer0_outputs(4329) <= inputs(218);
    layer0_outputs(4330) <= (inputs(192)) xor (inputs(91));
    layer0_outputs(4331) <= (inputs(212)) xor (inputs(180));
    layer0_outputs(4332) <= not(inputs(84)) or (inputs(14));
    layer0_outputs(4333) <= inputs(117);
    layer0_outputs(4334) <= inputs(176);
    layer0_outputs(4335) <= (inputs(116)) and not (inputs(211));
    layer0_outputs(4336) <= not(inputs(24));
    layer0_outputs(4337) <= (inputs(211)) and (inputs(245));
    layer0_outputs(4338) <= (inputs(110)) or (inputs(98));
    layer0_outputs(4339) <= not((inputs(243)) or (inputs(64)));
    layer0_outputs(4340) <= (inputs(115)) xor (inputs(254));
    layer0_outputs(4341) <= (inputs(61)) or (inputs(23));
    layer0_outputs(4342) <= inputs(38);
    layer0_outputs(4343) <= (inputs(97)) or (inputs(147));
    layer0_outputs(4344) <= (inputs(74)) or (inputs(170));
    layer0_outputs(4345) <= not(inputs(121));
    layer0_outputs(4346) <= (inputs(195)) or (inputs(62));
    layer0_outputs(4347) <= inputs(0);
    layer0_outputs(4348) <= not((inputs(238)) xor (inputs(250)));
    layer0_outputs(4349) <= (inputs(17)) and (inputs(79));
    layer0_outputs(4350) <= not(inputs(99)) or (inputs(188));
    layer0_outputs(4351) <= not(inputs(232));
    layer0_outputs(4352) <= (inputs(135)) or (inputs(31));
    layer0_outputs(4353) <= (inputs(126)) xor (inputs(207));
    layer0_outputs(4354) <= not((inputs(184)) or (inputs(133)));
    layer0_outputs(4355) <= '1';
    layer0_outputs(4356) <= not((inputs(77)) or (inputs(34)));
    layer0_outputs(4357) <= not(inputs(237));
    layer0_outputs(4358) <= (inputs(215)) and not (inputs(131));
    layer0_outputs(4359) <= (inputs(173)) and not (inputs(183));
    layer0_outputs(4360) <= (inputs(219)) or (inputs(155));
    layer0_outputs(4361) <= (inputs(15)) and not (inputs(192));
    layer0_outputs(4362) <= inputs(243);
    layer0_outputs(4363) <= not((inputs(70)) xor (inputs(99)));
    layer0_outputs(4364) <= not((inputs(168)) xor (inputs(15)));
    layer0_outputs(4365) <= inputs(138);
    layer0_outputs(4366) <= (inputs(66)) or (inputs(134));
    layer0_outputs(4367) <= not((inputs(43)) and (inputs(24)));
    layer0_outputs(4368) <= inputs(53);
    layer0_outputs(4369) <= inputs(232);
    layer0_outputs(4370) <= (inputs(153)) or (inputs(231));
    layer0_outputs(4371) <= (inputs(62)) and not (inputs(10));
    layer0_outputs(4372) <= (inputs(238)) xor (inputs(110));
    layer0_outputs(4373) <= (inputs(136)) and not (inputs(85));
    layer0_outputs(4374) <= (inputs(167)) or (inputs(212));
    layer0_outputs(4375) <= inputs(25);
    layer0_outputs(4376) <= not(inputs(102));
    layer0_outputs(4377) <= (inputs(112)) or (inputs(230));
    layer0_outputs(4378) <= not(inputs(243));
    layer0_outputs(4379) <= inputs(23);
    layer0_outputs(4380) <= not((inputs(79)) xor (inputs(230)));
    layer0_outputs(4381) <= not((inputs(232)) or (inputs(141)));
    layer0_outputs(4382) <= (inputs(111)) and (inputs(217));
    layer0_outputs(4383) <= inputs(228);
    layer0_outputs(4384) <= '0';
    layer0_outputs(4385) <= not(inputs(179));
    layer0_outputs(4386) <= (inputs(84)) and not (inputs(191));
    layer0_outputs(4387) <= (inputs(158)) or (inputs(75));
    layer0_outputs(4388) <= not(inputs(179)) or (inputs(244));
    layer0_outputs(4389) <= (inputs(125)) or (inputs(75));
    layer0_outputs(4390) <= not((inputs(225)) xor (inputs(199)));
    layer0_outputs(4391) <= (inputs(204)) or (inputs(107));
    layer0_outputs(4392) <= inputs(39);
    layer0_outputs(4393) <= inputs(106);
    layer0_outputs(4394) <= not(inputs(91));
    layer0_outputs(4395) <= not((inputs(198)) xor (inputs(242)));
    layer0_outputs(4396) <= not(inputs(126)) or (inputs(146));
    layer0_outputs(4397) <= (inputs(184)) and not (inputs(134));
    layer0_outputs(4398) <= not(inputs(118));
    layer0_outputs(4399) <= inputs(175);
    layer0_outputs(4400) <= not((inputs(63)) xor (inputs(143)));
    layer0_outputs(4401) <= not(inputs(139));
    layer0_outputs(4402) <= not((inputs(43)) or (inputs(97)));
    layer0_outputs(4403) <= '0';
    layer0_outputs(4404) <= not((inputs(206)) or (inputs(222)));
    layer0_outputs(4405) <= not(inputs(15)) or (inputs(95));
    layer0_outputs(4406) <= not(inputs(145)) or (inputs(117));
    layer0_outputs(4407) <= '1';
    layer0_outputs(4408) <= (inputs(208)) xor (inputs(165));
    layer0_outputs(4409) <= (inputs(76)) or (inputs(11));
    layer0_outputs(4410) <= (inputs(182)) and not (inputs(106));
    layer0_outputs(4411) <= not(inputs(216));
    layer0_outputs(4412) <= not((inputs(224)) and (inputs(204)));
    layer0_outputs(4413) <= not(inputs(149));
    layer0_outputs(4414) <= not((inputs(26)) and (inputs(65)));
    layer0_outputs(4415) <= inputs(81);
    layer0_outputs(4416) <= not((inputs(132)) or (inputs(20)));
    layer0_outputs(4417) <= '1';
    layer0_outputs(4418) <= not((inputs(78)) xor (inputs(156)));
    layer0_outputs(4419) <= not(inputs(228)) or (inputs(5));
    layer0_outputs(4420) <= (inputs(209)) or (inputs(202));
    layer0_outputs(4421) <= inputs(30);
    layer0_outputs(4422) <= not((inputs(20)) or (inputs(237)));
    layer0_outputs(4423) <= (inputs(111)) and (inputs(73));
    layer0_outputs(4424) <= not((inputs(176)) or (inputs(190)));
    layer0_outputs(4425) <= inputs(188);
    layer0_outputs(4426) <= not((inputs(83)) xor (inputs(54)));
    layer0_outputs(4427) <= (inputs(248)) and not (inputs(52));
    layer0_outputs(4428) <= not((inputs(176)) or (inputs(122)));
    layer0_outputs(4429) <= not(inputs(27));
    layer0_outputs(4430) <= '0';
    layer0_outputs(4431) <= (inputs(22)) xor (inputs(54));
    layer0_outputs(4432) <= (inputs(204)) and not (inputs(113));
    layer0_outputs(4433) <= (inputs(130)) and not (inputs(71));
    layer0_outputs(4434) <= not(inputs(126));
    layer0_outputs(4435) <= not((inputs(65)) xor (inputs(125)));
    layer0_outputs(4436) <= not(inputs(107)) or (inputs(160));
    layer0_outputs(4437) <= (inputs(138)) xor (inputs(198));
    layer0_outputs(4438) <= not((inputs(213)) or (inputs(82)));
    layer0_outputs(4439) <= not(inputs(147)) or (inputs(58));
    layer0_outputs(4440) <= not(inputs(202)) or (inputs(27));
    layer0_outputs(4441) <= not((inputs(253)) and (inputs(82)));
    layer0_outputs(4442) <= not(inputs(94));
    layer0_outputs(4443) <= not(inputs(83));
    layer0_outputs(4444) <= not((inputs(134)) xor (inputs(98)));
    layer0_outputs(4445) <= inputs(181);
    layer0_outputs(4446) <= inputs(157);
    layer0_outputs(4447) <= not(inputs(248));
    layer0_outputs(4448) <= not((inputs(15)) or (inputs(179)));
    layer0_outputs(4449) <= (inputs(71)) and not (inputs(197));
    layer0_outputs(4450) <= not(inputs(191)) or (inputs(142));
    layer0_outputs(4451) <= not(inputs(229)) or (inputs(139));
    layer0_outputs(4452) <= inputs(220);
    layer0_outputs(4453) <= (inputs(84)) xor (inputs(98));
    layer0_outputs(4454) <= not(inputs(29));
    layer0_outputs(4455) <= not(inputs(101)) or (inputs(103));
    layer0_outputs(4456) <= not(inputs(162));
    layer0_outputs(4457) <= (inputs(26)) or (inputs(238));
    layer0_outputs(4458) <= (inputs(169)) and (inputs(210));
    layer0_outputs(4459) <= not((inputs(210)) or (inputs(193)));
    layer0_outputs(4460) <= '0';
    layer0_outputs(4461) <= inputs(131);
    layer0_outputs(4462) <= (inputs(119)) and not (inputs(105));
    layer0_outputs(4463) <= (inputs(205)) or (inputs(184));
    layer0_outputs(4464) <= (inputs(135)) xor (inputs(34));
    layer0_outputs(4465) <= (inputs(110)) and not (inputs(135));
    layer0_outputs(4466) <= not((inputs(212)) and (inputs(185)));
    layer0_outputs(4467) <= '1';
    layer0_outputs(4468) <= inputs(29);
    layer0_outputs(4469) <= (inputs(143)) or (inputs(107));
    layer0_outputs(4470) <= not((inputs(104)) or (inputs(150)));
    layer0_outputs(4471) <= (inputs(9)) or (inputs(227));
    layer0_outputs(4472) <= (inputs(46)) or (inputs(117));
    layer0_outputs(4473) <= (inputs(203)) or (inputs(140));
    layer0_outputs(4474) <= not(inputs(249));
    layer0_outputs(4475) <= (inputs(200)) or (inputs(234));
    layer0_outputs(4476) <= inputs(196);
    layer0_outputs(4477) <= not((inputs(184)) or (inputs(94)));
    layer0_outputs(4478) <= not((inputs(195)) or (inputs(230)));
    layer0_outputs(4479) <= (inputs(105)) and not (inputs(150));
    layer0_outputs(4480) <= not((inputs(200)) and (inputs(207)));
    layer0_outputs(4481) <= (inputs(160)) xor (inputs(187));
    layer0_outputs(4482) <= (inputs(241)) and not (inputs(65));
    layer0_outputs(4483) <= inputs(71);
    layer0_outputs(4484) <= not((inputs(89)) xor (inputs(215)));
    layer0_outputs(4485) <= (inputs(252)) xor (inputs(134));
    layer0_outputs(4486) <= inputs(204);
    layer0_outputs(4487) <= not((inputs(44)) or (inputs(4)));
    layer0_outputs(4488) <= inputs(23);
    layer0_outputs(4489) <= not((inputs(142)) and (inputs(36)));
    layer0_outputs(4490) <= (inputs(155)) and not (inputs(29));
    layer0_outputs(4491) <= not((inputs(47)) or (inputs(42)));
    layer0_outputs(4492) <= '0';
    layer0_outputs(4493) <= (inputs(186)) xor (inputs(114));
    layer0_outputs(4494) <= (inputs(193)) xor (inputs(246));
    layer0_outputs(4495) <= not((inputs(177)) xor (inputs(47)));
    layer0_outputs(4496) <= (inputs(62)) and not (inputs(188));
    layer0_outputs(4497) <= inputs(165);
    layer0_outputs(4498) <= not(inputs(210));
    layer0_outputs(4499) <= (inputs(3)) or (inputs(192));
    layer0_outputs(4500) <= not((inputs(150)) or (inputs(58)));
    layer0_outputs(4501) <= inputs(104);
    layer0_outputs(4502) <= inputs(44);
    layer0_outputs(4503) <= not((inputs(8)) or (inputs(23)));
    layer0_outputs(4504) <= not((inputs(8)) xor (inputs(52)));
    layer0_outputs(4505) <= not(inputs(87)) or (inputs(143));
    layer0_outputs(4506) <= not((inputs(173)) xor (inputs(25)));
    layer0_outputs(4507) <= not(inputs(230));
    layer0_outputs(4508) <= (inputs(62)) and not (inputs(106));
    layer0_outputs(4509) <= (inputs(139)) or (inputs(174));
    layer0_outputs(4510) <= not(inputs(229));
    layer0_outputs(4511) <= not((inputs(107)) or (inputs(82)));
    layer0_outputs(4512) <= not(inputs(103));
    layer0_outputs(4513) <= (inputs(49)) xor (inputs(187));
    layer0_outputs(4514) <= not(inputs(84)) or (inputs(29));
    layer0_outputs(4515) <= '0';
    layer0_outputs(4516) <= (inputs(57)) and not (inputs(153));
    layer0_outputs(4517) <= (inputs(100)) and not (inputs(252));
    layer0_outputs(4518) <= not(inputs(198));
    layer0_outputs(4519) <= not((inputs(179)) or (inputs(70)));
    layer0_outputs(4520) <= (inputs(196)) or (inputs(187));
    layer0_outputs(4521) <= not((inputs(251)) and (inputs(65)));
    layer0_outputs(4522) <= inputs(232);
    layer0_outputs(4523) <= not(inputs(136)) or (inputs(4));
    layer0_outputs(4524) <= not(inputs(122)) or (inputs(16));
    layer0_outputs(4525) <= (inputs(95)) or (inputs(194));
    layer0_outputs(4526) <= not((inputs(122)) or (inputs(5)));
    layer0_outputs(4527) <= inputs(124);
    layer0_outputs(4528) <= inputs(120);
    layer0_outputs(4529) <= (inputs(27)) or (inputs(127));
    layer0_outputs(4530) <= not(inputs(83)) or (inputs(255));
    layer0_outputs(4531) <= not(inputs(165)) or (inputs(190));
    layer0_outputs(4532) <= not((inputs(245)) or (inputs(17)));
    layer0_outputs(4533) <= (inputs(173)) or (inputs(72));
    layer0_outputs(4534) <= inputs(171);
    layer0_outputs(4535) <= (inputs(32)) or (inputs(19));
    layer0_outputs(4536) <= (inputs(133)) and not (inputs(237));
    layer0_outputs(4537) <= not((inputs(74)) and (inputs(201)));
    layer0_outputs(4538) <= inputs(85);
    layer0_outputs(4539) <= not(inputs(87)) or (inputs(17));
    layer0_outputs(4540) <= not((inputs(96)) or (inputs(23)));
    layer0_outputs(4541) <= (inputs(17)) xor (inputs(41));
    layer0_outputs(4542) <= inputs(136);
    layer0_outputs(4543) <= (inputs(0)) or (inputs(33));
    layer0_outputs(4544) <= not((inputs(106)) xor (inputs(75)));
    layer0_outputs(4545) <= inputs(184);
    layer0_outputs(4546) <= not(inputs(249));
    layer0_outputs(4547) <= not(inputs(169));
    layer0_outputs(4548) <= (inputs(205)) and not (inputs(205));
    layer0_outputs(4549) <= (inputs(24)) and not (inputs(179));
    layer0_outputs(4550) <= not((inputs(72)) or (inputs(222)));
    layer0_outputs(4551) <= not(inputs(155));
    layer0_outputs(4552) <= not((inputs(182)) or (inputs(11)));
    layer0_outputs(4553) <= not(inputs(8)) or (inputs(12));
    layer0_outputs(4554) <= not(inputs(5)) or (inputs(158));
    layer0_outputs(4555) <= (inputs(189)) or (inputs(187));
    layer0_outputs(4556) <= (inputs(141)) and not (inputs(94));
    layer0_outputs(4557) <= not((inputs(142)) xor (inputs(75)));
    layer0_outputs(4558) <= not(inputs(200)) or (inputs(63));
    layer0_outputs(4559) <= (inputs(189)) or (inputs(220));
    layer0_outputs(4560) <= (inputs(166)) or (inputs(222));
    layer0_outputs(4561) <= (inputs(136)) and (inputs(60));
    layer0_outputs(4562) <= inputs(59);
    layer0_outputs(4563) <= not(inputs(179));
    layer0_outputs(4564) <= not(inputs(77));
    layer0_outputs(4565) <= not((inputs(19)) or (inputs(238)));
    layer0_outputs(4566) <= not((inputs(87)) and (inputs(77)));
    layer0_outputs(4567) <= not(inputs(228));
    layer0_outputs(4568) <= (inputs(243)) or (inputs(244));
    layer0_outputs(4569) <= (inputs(254)) or (inputs(2));
    layer0_outputs(4570) <= not((inputs(73)) and (inputs(111)));
    layer0_outputs(4571) <= (inputs(63)) xor (inputs(93));
    layer0_outputs(4572) <= '1';
    layer0_outputs(4573) <= not((inputs(255)) or (inputs(70)));
    layer0_outputs(4574) <= inputs(156);
    layer0_outputs(4575) <= not(inputs(39)) or (inputs(249));
    layer0_outputs(4576) <= not((inputs(185)) or (inputs(196)));
    layer0_outputs(4577) <= inputs(29);
    layer0_outputs(4578) <= not((inputs(143)) or (inputs(125)));
    layer0_outputs(4579) <= not(inputs(148));
    layer0_outputs(4580) <= not(inputs(78));
    layer0_outputs(4581) <= not((inputs(144)) or (inputs(163)));
    layer0_outputs(4582) <= (inputs(17)) or (inputs(193));
    layer0_outputs(4583) <= not(inputs(20)) or (inputs(248));
    layer0_outputs(4584) <= not(inputs(18)) or (inputs(247));
    layer0_outputs(4585) <= not(inputs(152));
    layer0_outputs(4586) <= inputs(175);
    layer0_outputs(4587) <= (inputs(192)) or (inputs(219));
    layer0_outputs(4588) <= (inputs(123)) and not (inputs(198));
    layer0_outputs(4589) <= not(inputs(215)) or (inputs(203));
    layer0_outputs(4590) <= (inputs(169)) or (inputs(223));
    layer0_outputs(4591) <= not(inputs(189));
    layer0_outputs(4592) <= inputs(184);
    layer0_outputs(4593) <= inputs(9);
    layer0_outputs(4594) <= inputs(181);
    layer0_outputs(4595) <= not(inputs(234)) or (inputs(178));
    layer0_outputs(4596) <= inputs(99);
    layer0_outputs(4597) <= (inputs(230)) xor (inputs(127));
    layer0_outputs(4598) <= inputs(136);
    layer0_outputs(4599) <= inputs(86);
    layer0_outputs(4600) <= (inputs(90)) xor (inputs(147));
    layer0_outputs(4601) <= inputs(110);
    layer0_outputs(4602) <= (inputs(208)) and not (inputs(47));
    layer0_outputs(4603) <= (inputs(67)) and not (inputs(238));
    layer0_outputs(4604) <= (inputs(157)) and not (inputs(238));
    layer0_outputs(4605) <= not((inputs(76)) xor (inputs(123)));
    layer0_outputs(4606) <= not((inputs(217)) or (inputs(144)));
    layer0_outputs(4607) <= not((inputs(226)) xor (inputs(127)));
    layer0_outputs(4608) <= not(inputs(228));
    layer0_outputs(4609) <= not(inputs(22));
    layer0_outputs(4610) <= not((inputs(64)) or (inputs(76)));
    layer0_outputs(4611) <= not(inputs(167));
    layer0_outputs(4612) <= not(inputs(177));
    layer0_outputs(4613) <= inputs(75);
    layer0_outputs(4614) <= not(inputs(189));
    layer0_outputs(4615) <= inputs(235);
    layer0_outputs(4616) <= (inputs(95)) xor (inputs(183));
    layer0_outputs(4617) <= inputs(200);
    layer0_outputs(4618) <= (inputs(57)) or (inputs(89));
    layer0_outputs(4619) <= inputs(93);
    layer0_outputs(4620) <= not((inputs(81)) xor (inputs(19)));
    layer0_outputs(4621) <= not((inputs(53)) xor (inputs(228)));
    layer0_outputs(4622) <= not(inputs(205));
    layer0_outputs(4623) <= inputs(97);
    layer0_outputs(4624) <= inputs(132);
    layer0_outputs(4625) <= not(inputs(161));
    layer0_outputs(4626) <= (inputs(231)) and not (inputs(79));
    layer0_outputs(4627) <= (inputs(187)) or (inputs(185));
    layer0_outputs(4628) <= (inputs(216)) and not (inputs(235));
    layer0_outputs(4629) <= not(inputs(138)) or (inputs(57));
    layer0_outputs(4630) <= (inputs(27)) or (inputs(113));
    layer0_outputs(4631) <= not(inputs(214)) or (inputs(5));
    layer0_outputs(4632) <= (inputs(103)) and not (inputs(61));
    layer0_outputs(4633) <= (inputs(1)) or (inputs(207));
    layer0_outputs(4634) <= not((inputs(228)) xor (inputs(239)));
    layer0_outputs(4635) <= not(inputs(113));
    layer0_outputs(4636) <= (inputs(234)) or (inputs(240));
    layer0_outputs(4637) <= (inputs(198)) or (inputs(184));
    layer0_outputs(4638) <= (inputs(238)) xor (inputs(59));
    layer0_outputs(4639) <= not(inputs(103));
    layer0_outputs(4640) <= inputs(136);
    layer0_outputs(4641) <= not((inputs(7)) or (inputs(67)));
    layer0_outputs(4642) <= inputs(86);
    layer0_outputs(4643) <= not((inputs(232)) xor (inputs(169)));
    layer0_outputs(4644) <= (inputs(195)) and not (inputs(67));
    layer0_outputs(4645) <= not(inputs(213)) or (inputs(92));
    layer0_outputs(4646) <= (inputs(57)) or (inputs(17));
    layer0_outputs(4647) <= not(inputs(231)) or (inputs(95));
    layer0_outputs(4648) <= not((inputs(212)) xor (inputs(149)));
    layer0_outputs(4649) <= (inputs(145)) xor (inputs(190));
    layer0_outputs(4650) <= inputs(211);
    layer0_outputs(4651) <= inputs(234);
    layer0_outputs(4652) <= '1';
    layer0_outputs(4653) <= '1';
    layer0_outputs(4654) <= (inputs(75)) and not (inputs(199));
    layer0_outputs(4655) <= not(inputs(163));
    layer0_outputs(4656) <= not((inputs(127)) or (inputs(63)));
    layer0_outputs(4657) <= not((inputs(210)) or (inputs(40)));
    layer0_outputs(4658) <= (inputs(218)) and not (inputs(248));
    layer0_outputs(4659) <= not(inputs(117));
    layer0_outputs(4660) <= not(inputs(93));
    layer0_outputs(4661) <= (inputs(141)) xor (inputs(205));
    layer0_outputs(4662) <= (inputs(114)) and not (inputs(247));
    layer0_outputs(4663) <= inputs(119);
    layer0_outputs(4664) <= '1';
    layer0_outputs(4665) <= not((inputs(238)) or (inputs(211)));
    layer0_outputs(4666) <= (inputs(139)) or (inputs(218));
    layer0_outputs(4667) <= (inputs(47)) or (inputs(115));
    layer0_outputs(4668) <= inputs(161);
    layer0_outputs(4669) <= (inputs(151)) or (inputs(240));
    layer0_outputs(4670) <= (inputs(230)) and (inputs(86));
    layer0_outputs(4671) <= '0';
    layer0_outputs(4672) <= not(inputs(164));
    layer0_outputs(4673) <= inputs(128);
    layer0_outputs(4674) <= (inputs(110)) or (inputs(2));
    layer0_outputs(4675) <= not(inputs(184));
    layer0_outputs(4676) <= (inputs(155)) xor (inputs(124));
    layer0_outputs(4677) <= not(inputs(43)) or (inputs(90));
    layer0_outputs(4678) <= inputs(209);
    layer0_outputs(4679) <= not(inputs(86));
    layer0_outputs(4680) <= not((inputs(85)) or (inputs(129)));
    layer0_outputs(4681) <= not((inputs(159)) and (inputs(58)));
    layer0_outputs(4682) <= not((inputs(196)) or (inputs(239)));
    layer0_outputs(4683) <= '0';
    layer0_outputs(4684) <= not((inputs(191)) or (inputs(227)));
    layer0_outputs(4685) <= inputs(105);
    layer0_outputs(4686) <= not(inputs(75));
    layer0_outputs(4687) <= not(inputs(54));
    layer0_outputs(4688) <= not((inputs(114)) xor (inputs(61)));
    layer0_outputs(4689) <= inputs(15);
    layer0_outputs(4690) <= (inputs(43)) and not (inputs(92));
    layer0_outputs(4691) <= (inputs(122)) or (inputs(125));
    layer0_outputs(4692) <= not(inputs(183)) or (inputs(68));
    layer0_outputs(4693) <= (inputs(224)) or (inputs(134));
    layer0_outputs(4694) <= not(inputs(78));
    layer0_outputs(4695) <= inputs(217);
    layer0_outputs(4696) <= inputs(198);
    layer0_outputs(4697) <= (inputs(21)) and not (inputs(170));
    layer0_outputs(4698) <= not((inputs(69)) xor (inputs(51)));
    layer0_outputs(4699) <= inputs(33);
    layer0_outputs(4700) <= (inputs(7)) or (inputs(84));
    layer0_outputs(4701) <= not((inputs(76)) or (inputs(126)));
    layer0_outputs(4702) <= (inputs(178)) or (inputs(69));
    layer0_outputs(4703) <= not(inputs(248));
    layer0_outputs(4704) <= (inputs(228)) and not (inputs(17));
    layer0_outputs(4705) <= inputs(54);
    layer0_outputs(4706) <= (inputs(166)) or (inputs(129));
    layer0_outputs(4707) <= (inputs(44)) and (inputs(61));
    layer0_outputs(4708) <= inputs(11);
    layer0_outputs(4709) <= not((inputs(228)) or (inputs(71)));
    layer0_outputs(4710) <= (inputs(59)) and (inputs(176));
    layer0_outputs(4711) <= not((inputs(229)) or (inputs(2)));
    layer0_outputs(4712) <= (inputs(176)) or (inputs(193));
    layer0_outputs(4713) <= not(inputs(48));
    layer0_outputs(4714) <= (inputs(88)) and not (inputs(1));
    layer0_outputs(4715) <= (inputs(109)) and not (inputs(236));
    layer0_outputs(4716) <= not((inputs(193)) xor (inputs(13)));
    layer0_outputs(4717) <= not(inputs(246));
    layer0_outputs(4718) <= (inputs(153)) or (inputs(64));
    layer0_outputs(4719) <= inputs(203);
    layer0_outputs(4720) <= (inputs(216)) and not (inputs(130));
    layer0_outputs(4721) <= not(inputs(114));
    layer0_outputs(4722) <= not((inputs(161)) xor (inputs(179)));
    layer0_outputs(4723) <= not(inputs(43));
    layer0_outputs(4724) <= not((inputs(251)) or (inputs(3)));
    layer0_outputs(4725) <= inputs(77);
    layer0_outputs(4726) <= (inputs(70)) xor (inputs(21));
    layer0_outputs(4727) <= (inputs(84)) xor (inputs(85));
    layer0_outputs(4728) <= (inputs(80)) and (inputs(121));
    layer0_outputs(4729) <= not(inputs(86)) or (inputs(92));
    layer0_outputs(4730) <= not(inputs(194)) or (inputs(47));
    layer0_outputs(4731) <= (inputs(11)) or (inputs(123));
    layer0_outputs(4732) <= (inputs(65)) and not (inputs(160));
    layer0_outputs(4733) <= not(inputs(253));
    layer0_outputs(4734) <= inputs(95);
    layer0_outputs(4735) <= inputs(165);
    layer0_outputs(4736) <= (inputs(82)) xor (inputs(201));
    layer0_outputs(4737) <= inputs(58);
    layer0_outputs(4738) <= not(inputs(225)) or (inputs(253));
    layer0_outputs(4739) <= (inputs(185)) and not (inputs(29));
    layer0_outputs(4740) <= '0';
    layer0_outputs(4741) <= inputs(178);
    layer0_outputs(4742) <= not((inputs(74)) and (inputs(149)));
    layer0_outputs(4743) <= not(inputs(101));
    layer0_outputs(4744) <= inputs(145);
    layer0_outputs(4745) <= not(inputs(140));
    layer0_outputs(4746) <= (inputs(116)) and not (inputs(173));
    layer0_outputs(4747) <= (inputs(181)) and not (inputs(95));
    layer0_outputs(4748) <= inputs(134);
    layer0_outputs(4749) <= not((inputs(29)) or (inputs(109)));
    layer0_outputs(4750) <= not(inputs(18));
    layer0_outputs(4751) <= inputs(136);
    layer0_outputs(4752) <= (inputs(180)) or (inputs(203));
    layer0_outputs(4753) <= not(inputs(168));
    layer0_outputs(4754) <= not(inputs(94)) or (inputs(236));
    layer0_outputs(4755) <= (inputs(219)) xor (inputs(24));
    layer0_outputs(4756) <= (inputs(139)) and (inputs(93));
    layer0_outputs(4757) <= inputs(231);
    layer0_outputs(4758) <= inputs(251);
    layer0_outputs(4759) <= not((inputs(14)) and (inputs(137)));
    layer0_outputs(4760) <= not(inputs(230));
    layer0_outputs(4761) <= not((inputs(135)) xor (inputs(128)));
    layer0_outputs(4762) <= not(inputs(238)) or (inputs(140));
    layer0_outputs(4763) <= not((inputs(234)) xor (inputs(225)));
    layer0_outputs(4764) <= not((inputs(189)) or (inputs(177)));
    layer0_outputs(4765) <= inputs(152);
    layer0_outputs(4766) <= (inputs(142)) or (inputs(218));
    layer0_outputs(4767) <= (inputs(121)) xor (inputs(193));
    layer0_outputs(4768) <= (inputs(121)) and not (inputs(132));
    layer0_outputs(4769) <= (inputs(16)) xor (inputs(61));
    layer0_outputs(4770) <= inputs(118);
    layer0_outputs(4771) <= not(inputs(45)) or (inputs(39));
    layer0_outputs(4772) <= not(inputs(42));
    layer0_outputs(4773) <= '1';
    layer0_outputs(4774) <= not(inputs(214));
    layer0_outputs(4775) <= inputs(179);
    layer0_outputs(4776) <= not((inputs(181)) or (inputs(187)));
    layer0_outputs(4777) <= (inputs(197)) and not (inputs(240));
    layer0_outputs(4778) <= not((inputs(44)) or (inputs(53)));
    layer0_outputs(4779) <= not(inputs(214)) or (inputs(81));
    layer0_outputs(4780) <= not((inputs(14)) or (inputs(5)));
    layer0_outputs(4781) <= inputs(224);
    layer0_outputs(4782) <= not(inputs(245));
    layer0_outputs(4783) <= not(inputs(33));
    layer0_outputs(4784) <= not(inputs(57)) or (inputs(249));
    layer0_outputs(4785) <= not(inputs(159)) or (inputs(4));
    layer0_outputs(4786) <= (inputs(71)) and not (inputs(191));
    layer0_outputs(4787) <= inputs(68);
    layer0_outputs(4788) <= not((inputs(231)) and (inputs(218)));
    layer0_outputs(4789) <= not(inputs(174)) or (inputs(184));
    layer0_outputs(4790) <= not(inputs(94)) or (inputs(15));
    layer0_outputs(4791) <= (inputs(54)) and not (inputs(91));
    layer0_outputs(4792) <= (inputs(42)) or (inputs(226));
    layer0_outputs(4793) <= (inputs(57)) and (inputs(50));
    layer0_outputs(4794) <= not((inputs(132)) or (inputs(56)));
    layer0_outputs(4795) <= inputs(232);
    layer0_outputs(4796) <= not(inputs(242)) or (inputs(127));
    layer0_outputs(4797) <= not((inputs(149)) or (inputs(237)));
    layer0_outputs(4798) <= (inputs(209)) or (inputs(160));
    layer0_outputs(4799) <= not((inputs(174)) or (inputs(135)));
    layer0_outputs(4800) <= (inputs(239)) and not (inputs(98));
    layer0_outputs(4801) <= not(inputs(104)) or (inputs(131));
    layer0_outputs(4802) <= not((inputs(60)) or (inputs(124)));
    layer0_outputs(4803) <= not(inputs(165));
    layer0_outputs(4804) <= not(inputs(246));
    layer0_outputs(4805) <= not((inputs(131)) xor (inputs(101)));
    layer0_outputs(4806) <= not(inputs(148)) or (inputs(183));
    layer0_outputs(4807) <= (inputs(92)) or (inputs(22));
    layer0_outputs(4808) <= not((inputs(153)) or (inputs(111)));
    layer0_outputs(4809) <= '1';
    layer0_outputs(4810) <= (inputs(161)) and not (inputs(59));
    layer0_outputs(4811) <= (inputs(3)) or (inputs(219));
    layer0_outputs(4812) <= not(inputs(247)) or (inputs(79));
    layer0_outputs(4813) <= not(inputs(243));
    layer0_outputs(4814) <= not(inputs(224));
    layer0_outputs(4815) <= '0';
    layer0_outputs(4816) <= not(inputs(104));
    layer0_outputs(4817) <= not(inputs(208));
    layer0_outputs(4818) <= (inputs(26)) or (inputs(97));
    layer0_outputs(4819) <= (inputs(97)) and not (inputs(73));
    layer0_outputs(4820) <= (inputs(228)) or (inputs(246));
    layer0_outputs(4821) <= (inputs(199)) xor (inputs(214));
    layer0_outputs(4822) <= '0';
    layer0_outputs(4823) <= not((inputs(160)) xor (inputs(24)));
    layer0_outputs(4824) <= not(inputs(7)) or (inputs(191));
    layer0_outputs(4825) <= inputs(53);
    layer0_outputs(4826) <= not(inputs(157)) or (inputs(239));
    layer0_outputs(4827) <= inputs(178);
    layer0_outputs(4828) <= (inputs(66)) and not (inputs(182));
    layer0_outputs(4829) <= not(inputs(198)) or (inputs(133));
    layer0_outputs(4830) <= '0';
    layer0_outputs(4831) <= not(inputs(168)) or (inputs(118));
    layer0_outputs(4832) <= not(inputs(76));
    layer0_outputs(4833) <= (inputs(206)) or (inputs(168));
    layer0_outputs(4834) <= not(inputs(222)) or (inputs(72));
    layer0_outputs(4835) <= inputs(156);
    layer0_outputs(4836) <= (inputs(247)) and not (inputs(236));
    layer0_outputs(4837) <= not(inputs(156));
    layer0_outputs(4838) <= inputs(24);
    layer0_outputs(4839) <= not((inputs(136)) or (inputs(192)));
    layer0_outputs(4840) <= not((inputs(171)) xor (inputs(172)));
    layer0_outputs(4841) <= inputs(60);
    layer0_outputs(4842) <= (inputs(121)) and not (inputs(180));
    layer0_outputs(4843) <= (inputs(193)) and not (inputs(109));
    layer0_outputs(4844) <= (inputs(54)) or (inputs(109));
    layer0_outputs(4845) <= not((inputs(79)) xor (inputs(12)));
    layer0_outputs(4846) <= inputs(20);
    layer0_outputs(4847) <= inputs(60);
    layer0_outputs(4848) <= not(inputs(73));
    layer0_outputs(4849) <= '0';
    layer0_outputs(4850) <= not((inputs(93)) or (inputs(188)));
    layer0_outputs(4851) <= inputs(124);
    layer0_outputs(4852) <= not(inputs(169)) or (inputs(144));
    layer0_outputs(4853) <= '0';
    layer0_outputs(4854) <= not(inputs(124));
    layer0_outputs(4855) <= not((inputs(185)) or (inputs(49)));
    layer0_outputs(4856) <= inputs(84);
    layer0_outputs(4857) <= (inputs(253)) or (inputs(231));
    layer0_outputs(4858) <= not(inputs(119));
    layer0_outputs(4859) <= (inputs(195)) or (inputs(223));
    layer0_outputs(4860) <= (inputs(222)) or (inputs(32));
    layer0_outputs(4861) <= not((inputs(251)) xor (inputs(2)));
    layer0_outputs(4862) <= '1';
    layer0_outputs(4863) <= inputs(227);
    layer0_outputs(4864) <= not(inputs(126)) or (inputs(78));
    layer0_outputs(4865) <= (inputs(244)) or (inputs(209));
    layer0_outputs(4866) <= not((inputs(18)) xor (inputs(81)));
    layer0_outputs(4867) <= not(inputs(159));
    layer0_outputs(4868) <= not(inputs(39)) or (inputs(198));
    layer0_outputs(4869) <= not((inputs(207)) or (inputs(39)));
    layer0_outputs(4870) <= not(inputs(10));
    layer0_outputs(4871) <= (inputs(194)) and not (inputs(175));
    layer0_outputs(4872) <= inputs(235);
    layer0_outputs(4873) <= not((inputs(246)) and (inputs(28)));
    layer0_outputs(4874) <= not((inputs(86)) xor (inputs(225)));
    layer0_outputs(4875) <= not(inputs(88)) or (inputs(15));
    layer0_outputs(4876) <= not(inputs(0));
    layer0_outputs(4877) <= inputs(195);
    layer0_outputs(4878) <= (inputs(213)) or (inputs(3));
    layer0_outputs(4879) <= (inputs(56)) and (inputs(59));
    layer0_outputs(4880) <= inputs(130);
    layer0_outputs(4881) <= inputs(109);
    layer0_outputs(4882) <= inputs(210);
    layer0_outputs(4883) <= inputs(134);
    layer0_outputs(4884) <= not(inputs(121));
    layer0_outputs(4885) <= '1';
    layer0_outputs(4886) <= (inputs(43)) or (inputs(97));
    layer0_outputs(4887) <= inputs(7);
    layer0_outputs(4888) <= inputs(69);
    layer0_outputs(4889) <= not(inputs(46));
    layer0_outputs(4890) <= not((inputs(205)) or (inputs(145)));
    layer0_outputs(4891) <= (inputs(45)) xor (inputs(76));
    layer0_outputs(4892) <= (inputs(107)) and not (inputs(87));
    layer0_outputs(4893) <= not(inputs(149));
    layer0_outputs(4894) <= not(inputs(180)) or (inputs(0));
    layer0_outputs(4895) <= inputs(23);
    layer0_outputs(4896) <= not(inputs(76)) or (inputs(171));
    layer0_outputs(4897) <= not(inputs(72));
    layer0_outputs(4898) <= (inputs(46)) or (inputs(197));
    layer0_outputs(4899) <= (inputs(8)) or (inputs(62));
    layer0_outputs(4900) <= not((inputs(84)) xor (inputs(192)));
    layer0_outputs(4901) <= not((inputs(31)) xor (inputs(116)));
    layer0_outputs(4902) <= inputs(125);
    layer0_outputs(4903) <= (inputs(171)) xor (inputs(205));
    layer0_outputs(4904) <= (inputs(23)) and not (inputs(234));
    layer0_outputs(4905) <= (inputs(196)) and not (inputs(221));
    layer0_outputs(4906) <= (inputs(172)) and (inputs(57));
    layer0_outputs(4907) <= inputs(180);
    layer0_outputs(4908) <= (inputs(147)) and not (inputs(14));
    layer0_outputs(4909) <= not((inputs(68)) or (inputs(197)));
    layer0_outputs(4910) <= not(inputs(233)) or (inputs(52));
    layer0_outputs(4911) <= not((inputs(34)) or (inputs(2)));
    layer0_outputs(4912) <= not(inputs(80)) or (inputs(199));
    layer0_outputs(4913) <= not(inputs(97));
    layer0_outputs(4914) <= not((inputs(15)) or (inputs(169)));
    layer0_outputs(4915) <= (inputs(182)) or (inputs(254));
    layer0_outputs(4916) <= not((inputs(156)) or (inputs(59)));
    layer0_outputs(4917) <= (inputs(87)) or (inputs(81));
    layer0_outputs(4918) <= not(inputs(105));
    layer0_outputs(4919) <= inputs(234);
    layer0_outputs(4920) <= inputs(167);
    layer0_outputs(4921) <= not(inputs(151));
    layer0_outputs(4922) <= not(inputs(107)) or (inputs(183));
    layer0_outputs(4923) <= not(inputs(175));
    layer0_outputs(4924) <= inputs(159);
    layer0_outputs(4925) <= (inputs(160)) and not (inputs(15));
    layer0_outputs(4926) <= not(inputs(99));
    layer0_outputs(4927) <= not((inputs(116)) or (inputs(97)));
    layer0_outputs(4928) <= not((inputs(108)) or (inputs(254)));
    layer0_outputs(4929) <= not(inputs(27)) or (inputs(116));
    layer0_outputs(4930) <= (inputs(186)) or (inputs(252));
    layer0_outputs(4931) <= inputs(3);
    layer0_outputs(4932) <= (inputs(187)) and not (inputs(4));
    layer0_outputs(4933) <= (inputs(4)) and not (inputs(157));
    layer0_outputs(4934) <= inputs(232);
    layer0_outputs(4935) <= inputs(220);
    layer0_outputs(4936) <= inputs(160);
    layer0_outputs(4937) <= inputs(217);
    layer0_outputs(4938) <= not(inputs(219));
    layer0_outputs(4939) <= not((inputs(208)) xor (inputs(22)));
    layer0_outputs(4940) <= (inputs(243)) or (inputs(125));
    layer0_outputs(4941) <= not(inputs(217)) or (inputs(59));
    layer0_outputs(4942) <= not(inputs(40));
    layer0_outputs(4943) <= not((inputs(178)) or (inputs(179)));
    layer0_outputs(4944) <= (inputs(139)) xor (inputs(118));
    layer0_outputs(4945) <= inputs(120);
    layer0_outputs(4946) <= not((inputs(179)) or (inputs(212)));
    layer0_outputs(4947) <= '1';
    layer0_outputs(4948) <= not((inputs(178)) xor (inputs(82)));
    layer0_outputs(4949) <= inputs(234);
    layer0_outputs(4950) <= inputs(60);
    layer0_outputs(4951) <= not(inputs(90));
    layer0_outputs(4952) <= (inputs(139)) or (inputs(12));
    layer0_outputs(4953) <= '1';
    layer0_outputs(4954) <= not(inputs(240));
    layer0_outputs(4955) <= not(inputs(91));
    layer0_outputs(4956) <= inputs(26);
    layer0_outputs(4957) <= inputs(150);
    layer0_outputs(4958) <= not((inputs(46)) or (inputs(243)));
    layer0_outputs(4959) <= (inputs(21)) and not (inputs(129));
    layer0_outputs(4960) <= (inputs(82)) and not (inputs(88));
    layer0_outputs(4961) <= not(inputs(233));
    layer0_outputs(4962) <= not((inputs(244)) or (inputs(220)));
    layer0_outputs(4963) <= (inputs(1)) or (inputs(197));
    layer0_outputs(4964) <= not(inputs(154));
    layer0_outputs(4965) <= (inputs(123)) and (inputs(108));
    layer0_outputs(4966) <= (inputs(119)) or (inputs(183));
    layer0_outputs(4967) <= not((inputs(102)) xor (inputs(158)));
    layer0_outputs(4968) <= not(inputs(219)) or (inputs(246));
    layer0_outputs(4969) <= not(inputs(130));
    layer0_outputs(4970) <= inputs(30);
    layer0_outputs(4971) <= (inputs(175)) xor (inputs(78));
    layer0_outputs(4972) <= '1';
    layer0_outputs(4973) <= (inputs(218)) and not (inputs(67));
    layer0_outputs(4974) <= inputs(88);
    layer0_outputs(4975) <= (inputs(26)) or (inputs(63));
    layer0_outputs(4976) <= (inputs(84)) or (inputs(160));
    layer0_outputs(4977) <= not(inputs(190)) or (inputs(197));
    layer0_outputs(4978) <= not(inputs(190)) or (inputs(120));
    layer0_outputs(4979) <= not(inputs(113));
    layer0_outputs(4980) <= inputs(81);
    layer0_outputs(4981) <= (inputs(190)) or (inputs(153));
    layer0_outputs(4982) <= not(inputs(104)) or (inputs(97));
    layer0_outputs(4983) <= inputs(44);
    layer0_outputs(4984) <= inputs(174);
    layer0_outputs(4985) <= not((inputs(167)) xor (inputs(164)));
    layer0_outputs(4986) <= '1';
    layer0_outputs(4987) <= (inputs(109)) or (inputs(162));
    layer0_outputs(4988) <= not(inputs(15));
    layer0_outputs(4989) <= (inputs(245)) and not (inputs(165));
    layer0_outputs(4990) <= not(inputs(252)) or (inputs(47));
    layer0_outputs(4991) <= not(inputs(206)) or (inputs(40));
    layer0_outputs(4992) <= not((inputs(188)) and (inputs(200)));
    layer0_outputs(4993) <= inputs(78);
    layer0_outputs(4994) <= not(inputs(179));
    layer0_outputs(4995) <= (inputs(163)) or (inputs(126));
    layer0_outputs(4996) <= not((inputs(77)) or (inputs(169)));
    layer0_outputs(4997) <= (inputs(18)) and not (inputs(51));
    layer0_outputs(4998) <= not(inputs(209)) or (inputs(87));
    layer0_outputs(4999) <= (inputs(229)) and not (inputs(166));
    layer0_outputs(5000) <= not((inputs(172)) xor (inputs(236)));
    layer0_outputs(5001) <= (inputs(64)) or (inputs(56));
    layer0_outputs(5002) <= not(inputs(113));
    layer0_outputs(5003) <= not((inputs(201)) and (inputs(211)));
    layer0_outputs(5004) <= not((inputs(222)) or (inputs(110)));
    layer0_outputs(5005) <= not(inputs(173));
    layer0_outputs(5006) <= not(inputs(49));
    layer0_outputs(5007) <= inputs(161);
    layer0_outputs(5008) <= not(inputs(201)) or (inputs(110));
    layer0_outputs(5009) <= (inputs(222)) and (inputs(226));
    layer0_outputs(5010) <= not(inputs(100)) or (inputs(168));
    layer0_outputs(5011) <= not((inputs(185)) or (inputs(104)));
    layer0_outputs(5012) <= not(inputs(116));
    layer0_outputs(5013) <= not(inputs(36)) or (inputs(8));
    layer0_outputs(5014) <= (inputs(191)) or (inputs(53));
    layer0_outputs(5015) <= not(inputs(78));
    layer0_outputs(5016) <= (inputs(1)) or (inputs(128));
    layer0_outputs(5017) <= not(inputs(120));
    layer0_outputs(5018) <= (inputs(204)) or (inputs(236));
    layer0_outputs(5019) <= not(inputs(247));
    layer0_outputs(5020) <= not((inputs(238)) or (inputs(221)));
    layer0_outputs(5021) <= not(inputs(159)) or (inputs(16));
    layer0_outputs(5022) <= not(inputs(69)) or (inputs(255));
    layer0_outputs(5023) <= (inputs(78)) and (inputs(182));
    layer0_outputs(5024) <= not((inputs(203)) xor (inputs(231)));
    layer0_outputs(5025) <= (inputs(95)) or (inputs(210));
    layer0_outputs(5026) <= (inputs(137)) and not (inputs(18));
    layer0_outputs(5027) <= inputs(37);
    layer0_outputs(5028) <= not((inputs(142)) or (inputs(10)));
    layer0_outputs(5029) <= not(inputs(163)) or (inputs(11));
    layer0_outputs(5030) <= not((inputs(38)) or (inputs(146)));
    layer0_outputs(5031) <= (inputs(218)) and (inputs(131));
    layer0_outputs(5032) <= (inputs(88)) or (inputs(241));
    layer0_outputs(5033) <= (inputs(97)) and (inputs(177));
    layer0_outputs(5034) <= not(inputs(208));
    layer0_outputs(5035) <= (inputs(208)) or (inputs(254));
    layer0_outputs(5036) <= inputs(140);
    layer0_outputs(5037) <= not(inputs(205)) or (inputs(255));
    layer0_outputs(5038) <= (inputs(185)) and not (inputs(100));
    layer0_outputs(5039) <= not((inputs(111)) or (inputs(172)));
    layer0_outputs(5040) <= not(inputs(75)) or (inputs(7));
    layer0_outputs(5041) <= not((inputs(73)) or (inputs(117)));
    layer0_outputs(5042) <= (inputs(252)) and (inputs(51));
    layer0_outputs(5043) <= '0';
    layer0_outputs(5044) <= inputs(29);
    layer0_outputs(5045) <= (inputs(44)) xor (inputs(3));
    layer0_outputs(5046) <= not(inputs(135));
    layer0_outputs(5047) <= inputs(251);
    layer0_outputs(5048) <= (inputs(161)) or (inputs(147));
    layer0_outputs(5049) <= not(inputs(229)) or (inputs(81));
    layer0_outputs(5050) <= (inputs(34)) or (inputs(60));
    layer0_outputs(5051) <= not(inputs(118));
    layer0_outputs(5052) <= inputs(112);
    layer0_outputs(5053) <= (inputs(159)) or (inputs(193));
    layer0_outputs(5054) <= not(inputs(104));
    layer0_outputs(5055) <= (inputs(211)) or (inputs(80));
    layer0_outputs(5056) <= not((inputs(155)) xor (inputs(197)));
    layer0_outputs(5057) <= not((inputs(167)) or (inputs(191)));
    layer0_outputs(5058) <= not(inputs(185));
    layer0_outputs(5059) <= (inputs(187)) and not (inputs(239));
    layer0_outputs(5060) <= not(inputs(166));
    layer0_outputs(5061) <= inputs(194);
    layer0_outputs(5062) <= (inputs(31)) or (inputs(178));
    layer0_outputs(5063) <= inputs(206);
    layer0_outputs(5064) <= not(inputs(160)) or (inputs(105));
    layer0_outputs(5065) <= (inputs(70)) and not (inputs(76));
    layer0_outputs(5066) <= not((inputs(172)) and (inputs(232)));
    layer0_outputs(5067) <= not(inputs(89)) or (inputs(33));
    layer0_outputs(5068) <= (inputs(90)) xor (inputs(21));
    layer0_outputs(5069) <= (inputs(56)) and not (inputs(133));
    layer0_outputs(5070) <= (inputs(128)) and not (inputs(255));
    layer0_outputs(5071) <= inputs(110);
    layer0_outputs(5072) <= (inputs(0)) or (inputs(246));
    layer0_outputs(5073) <= (inputs(194)) or (inputs(235));
    layer0_outputs(5074) <= not(inputs(170));
    layer0_outputs(5075) <= (inputs(188)) or (inputs(236));
    layer0_outputs(5076) <= (inputs(103)) and not (inputs(166));
    layer0_outputs(5077) <= not(inputs(213));
    layer0_outputs(5078) <= (inputs(122)) and not (inputs(255));
    layer0_outputs(5079) <= not(inputs(140));
    layer0_outputs(5080) <= not(inputs(75)) or (inputs(40));
    layer0_outputs(5081) <= inputs(152);
    layer0_outputs(5082) <= inputs(206);
    layer0_outputs(5083) <= not(inputs(246)) or (inputs(33));
    layer0_outputs(5084) <= not((inputs(202)) xor (inputs(89)));
    layer0_outputs(5085) <= (inputs(156)) xor (inputs(33));
    layer0_outputs(5086) <= not(inputs(107)) or (inputs(219));
    layer0_outputs(5087) <= not(inputs(43));
    layer0_outputs(5088) <= (inputs(204)) and not (inputs(63));
    layer0_outputs(5089) <= (inputs(81)) or (inputs(236));
    layer0_outputs(5090) <= not(inputs(228));
    layer0_outputs(5091) <= (inputs(38)) or (inputs(114));
    layer0_outputs(5092) <= (inputs(17)) and not (inputs(77));
    layer0_outputs(5093) <= inputs(92);
    layer0_outputs(5094) <= (inputs(84)) or (inputs(50));
    layer0_outputs(5095) <= not(inputs(163));
    layer0_outputs(5096) <= inputs(234);
    layer0_outputs(5097) <= not((inputs(181)) xor (inputs(59)));
    layer0_outputs(5098) <= not(inputs(227));
    layer0_outputs(5099) <= not(inputs(97));
    layer0_outputs(5100) <= (inputs(217)) and (inputs(133));
    layer0_outputs(5101) <= not((inputs(187)) or (inputs(20)));
    layer0_outputs(5102) <= (inputs(53)) xor (inputs(223));
    layer0_outputs(5103) <= (inputs(46)) xor (inputs(4));
    layer0_outputs(5104) <= not((inputs(96)) xor (inputs(26)));
    layer0_outputs(5105) <= (inputs(24)) and (inputs(42));
    layer0_outputs(5106) <= not(inputs(132));
    layer0_outputs(5107) <= (inputs(192)) or (inputs(214));
    layer0_outputs(5108) <= (inputs(200)) and (inputs(96));
    layer0_outputs(5109) <= inputs(20);
    layer0_outputs(5110) <= not((inputs(85)) xor (inputs(102)));
    layer0_outputs(5111) <= (inputs(141)) and (inputs(226));
    layer0_outputs(5112) <= not((inputs(111)) or (inputs(93)));
    layer0_outputs(5113) <= (inputs(198)) or (inputs(174));
    layer0_outputs(5114) <= inputs(219);
    layer0_outputs(5115) <= (inputs(39)) xor (inputs(52));
    layer0_outputs(5116) <= inputs(41);
    layer0_outputs(5117) <= not(inputs(203)) or (inputs(153));
    layer0_outputs(5118) <= (inputs(231)) and (inputs(131));
    layer0_outputs(5119) <= not(inputs(246)) or (inputs(95));
    layer0_outputs(5120) <= not((inputs(105)) or (inputs(76)));
    layer0_outputs(5121) <= not(inputs(146));
    layer0_outputs(5122) <= not((inputs(181)) or (inputs(92)));
    layer0_outputs(5123) <= not((inputs(231)) and (inputs(42)));
    layer0_outputs(5124) <= not(inputs(111));
    layer0_outputs(5125) <= '1';
    layer0_outputs(5126) <= not(inputs(23));
    layer0_outputs(5127) <= (inputs(56)) and not (inputs(148));
    layer0_outputs(5128) <= not(inputs(119));
    layer0_outputs(5129) <= (inputs(137)) xor (inputs(142));
    layer0_outputs(5130) <= (inputs(145)) and (inputs(143));
    layer0_outputs(5131) <= not(inputs(163));
    layer0_outputs(5132) <= (inputs(250)) and not (inputs(98));
    layer0_outputs(5133) <= (inputs(83)) and not (inputs(143));
    layer0_outputs(5134) <= (inputs(130)) xor (inputs(148));
    layer0_outputs(5135) <= inputs(245);
    layer0_outputs(5136) <= not((inputs(63)) xor (inputs(143)));
    layer0_outputs(5137) <= not(inputs(184));
    layer0_outputs(5138) <= not(inputs(152)) or (inputs(47));
    layer0_outputs(5139) <= not(inputs(244));
    layer0_outputs(5140) <= not(inputs(173)) or (inputs(112));
    layer0_outputs(5141) <= not(inputs(26));
    layer0_outputs(5142) <= inputs(231);
    layer0_outputs(5143) <= not((inputs(134)) or (inputs(198)));
    layer0_outputs(5144) <= (inputs(44)) and (inputs(186));
    layer0_outputs(5145) <= not(inputs(230));
    layer0_outputs(5146) <= (inputs(57)) and (inputs(117));
    layer0_outputs(5147) <= (inputs(76)) or (inputs(53));
    layer0_outputs(5148) <= (inputs(72)) xor (inputs(60));
    layer0_outputs(5149) <= inputs(102);
    layer0_outputs(5150) <= not(inputs(65));
    layer0_outputs(5151) <= not(inputs(193));
    layer0_outputs(5152) <= not(inputs(101)) or (inputs(66));
    layer0_outputs(5153) <= not(inputs(28)) or (inputs(5));
    layer0_outputs(5154) <= (inputs(205)) or (inputs(250));
    layer0_outputs(5155) <= (inputs(42)) and (inputs(211));
    layer0_outputs(5156) <= not(inputs(60)) or (inputs(183));
    layer0_outputs(5157) <= (inputs(131)) or (inputs(211));
    layer0_outputs(5158) <= not(inputs(54)) or (inputs(154));
    layer0_outputs(5159) <= (inputs(124)) and not (inputs(161));
    layer0_outputs(5160) <= inputs(69);
    layer0_outputs(5161) <= not((inputs(80)) or (inputs(226)));
    layer0_outputs(5162) <= (inputs(168)) and not (inputs(30));
    layer0_outputs(5163) <= not(inputs(64)) or (inputs(44));
    layer0_outputs(5164) <= not(inputs(99));
    layer0_outputs(5165) <= '1';
    layer0_outputs(5166) <= not(inputs(105));
    layer0_outputs(5167) <= not((inputs(140)) and (inputs(254)));
    layer0_outputs(5168) <= not(inputs(75)) or (inputs(35));
    layer0_outputs(5169) <= (inputs(100)) and not (inputs(193));
    layer0_outputs(5170) <= (inputs(72)) or (inputs(209));
    layer0_outputs(5171) <= not((inputs(44)) or (inputs(91)));
    layer0_outputs(5172) <= (inputs(167)) or (inputs(103));
    layer0_outputs(5173) <= inputs(86);
    layer0_outputs(5174) <= not((inputs(205)) or (inputs(227)));
    layer0_outputs(5175) <= not(inputs(45)) or (inputs(226));
    layer0_outputs(5176) <= (inputs(162)) or (inputs(98));
    layer0_outputs(5177) <= (inputs(71)) and not (inputs(13));
    layer0_outputs(5178) <= not(inputs(25));
    layer0_outputs(5179) <= not(inputs(42));
    layer0_outputs(5180) <= not((inputs(111)) or (inputs(174)));
    layer0_outputs(5181) <= not(inputs(122)) or (inputs(176));
    layer0_outputs(5182) <= not((inputs(166)) or (inputs(104)));
    layer0_outputs(5183) <= not((inputs(195)) or (inputs(162)));
    layer0_outputs(5184) <= (inputs(226)) and not (inputs(152));
    layer0_outputs(5185) <= not(inputs(29));
    layer0_outputs(5186) <= '1';
    layer0_outputs(5187) <= not(inputs(10)) or (inputs(82));
    layer0_outputs(5188) <= (inputs(202)) and (inputs(216));
    layer0_outputs(5189) <= inputs(134);
    layer0_outputs(5190) <= '1';
    layer0_outputs(5191) <= '0';
    layer0_outputs(5192) <= inputs(113);
    layer0_outputs(5193) <= not((inputs(73)) or (inputs(240)));
    layer0_outputs(5194) <= not(inputs(246));
    layer0_outputs(5195) <= '1';
    layer0_outputs(5196) <= (inputs(71)) or (inputs(250));
    layer0_outputs(5197) <= not((inputs(22)) and (inputs(40)));
    layer0_outputs(5198) <= not(inputs(178)) or (inputs(163));
    layer0_outputs(5199) <= not(inputs(191)) or (inputs(29));
    layer0_outputs(5200) <= not((inputs(213)) or (inputs(144)));
    layer0_outputs(5201) <= (inputs(118)) and not (inputs(237));
    layer0_outputs(5202) <= (inputs(50)) xor (inputs(108));
    layer0_outputs(5203) <= not(inputs(65)) or (inputs(250));
    layer0_outputs(5204) <= not((inputs(245)) xor (inputs(244)));
    layer0_outputs(5205) <= not((inputs(207)) or (inputs(192)));
    layer0_outputs(5206) <= not(inputs(35)) or (inputs(75));
    layer0_outputs(5207) <= not(inputs(85));
    layer0_outputs(5208) <= (inputs(231)) and not (inputs(75));
    layer0_outputs(5209) <= (inputs(233)) xor (inputs(207));
    layer0_outputs(5210) <= (inputs(7)) and not (inputs(161));
    layer0_outputs(5211) <= not(inputs(126));
    layer0_outputs(5212) <= inputs(132);
    layer0_outputs(5213) <= not(inputs(25)) or (inputs(179));
    layer0_outputs(5214) <= (inputs(71)) xor (inputs(27));
    layer0_outputs(5215) <= (inputs(68)) and not (inputs(245));
    layer0_outputs(5216) <= inputs(18);
    layer0_outputs(5217) <= not((inputs(55)) and (inputs(193)));
    layer0_outputs(5218) <= not((inputs(196)) xor (inputs(179)));
    layer0_outputs(5219) <= (inputs(7)) or (inputs(203));
    layer0_outputs(5220) <= not((inputs(202)) or (inputs(222)));
    layer0_outputs(5221) <= not(inputs(110)) or (inputs(35));
    layer0_outputs(5222) <= (inputs(199)) and (inputs(58));
    layer0_outputs(5223) <= inputs(104);
    layer0_outputs(5224) <= not((inputs(67)) or (inputs(49)));
    layer0_outputs(5225) <= not(inputs(110)) or (inputs(223));
    layer0_outputs(5226) <= (inputs(184)) and not (inputs(71));
    layer0_outputs(5227) <= inputs(95);
    layer0_outputs(5228) <= not(inputs(95)) or (inputs(88));
    layer0_outputs(5229) <= (inputs(232)) or (inputs(251));
    layer0_outputs(5230) <= not(inputs(103)) or (inputs(125));
    layer0_outputs(5231) <= inputs(42);
    layer0_outputs(5232) <= not(inputs(100)) or (inputs(215));
    layer0_outputs(5233) <= inputs(135);
    layer0_outputs(5234) <= inputs(89);
    layer0_outputs(5235) <= inputs(152);
    layer0_outputs(5236) <= inputs(150);
    layer0_outputs(5237) <= not((inputs(128)) and (inputs(160)));
    layer0_outputs(5238) <= not((inputs(7)) xor (inputs(95)));
    layer0_outputs(5239) <= inputs(152);
    layer0_outputs(5240) <= not(inputs(134)) or (inputs(238));
    layer0_outputs(5241) <= not(inputs(247));
    layer0_outputs(5242) <= inputs(167);
    layer0_outputs(5243) <= not(inputs(116));
    layer0_outputs(5244) <= inputs(117);
    layer0_outputs(5245) <= not((inputs(146)) or (inputs(113)));
    layer0_outputs(5246) <= not((inputs(133)) or (inputs(40)));
    layer0_outputs(5247) <= (inputs(22)) xor (inputs(236));
    layer0_outputs(5248) <= '1';
    layer0_outputs(5249) <= not(inputs(141));
    layer0_outputs(5250) <= inputs(243);
    layer0_outputs(5251) <= (inputs(214)) and not (inputs(38));
    layer0_outputs(5252) <= not((inputs(132)) and (inputs(116)));
    layer0_outputs(5253) <= (inputs(68)) xor (inputs(232));
    layer0_outputs(5254) <= not(inputs(242)) or (inputs(47));
    layer0_outputs(5255) <= not((inputs(1)) xor (inputs(130)));
    layer0_outputs(5256) <= (inputs(189)) and not (inputs(88));
    layer0_outputs(5257) <= not(inputs(155)) or (inputs(237));
    layer0_outputs(5258) <= inputs(204);
    layer0_outputs(5259) <= (inputs(219)) and (inputs(240));
    layer0_outputs(5260) <= (inputs(100)) xor (inputs(65));
    layer0_outputs(5261) <= not(inputs(14)) or (inputs(198));
    layer0_outputs(5262) <= (inputs(122)) or (inputs(78));
    layer0_outputs(5263) <= inputs(86);
    layer0_outputs(5264) <= not((inputs(86)) or (inputs(68)));
    layer0_outputs(5265) <= not((inputs(9)) xor (inputs(41)));
    layer0_outputs(5266) <= (inputs(240)) and not (inputs(65));
    layer0_outputs(5267) <= inputs(143);
    layer0_outputs(5268) <= (inputs(223)) or (inputs(188));
    layer0_outputs(5269) <= inputs(182);
    layer0_outputs(5270) <= not(inputs(25));
    layer0_outputs(5271) <= (inputs(117)) or (inputs(84));
    layer0_outputs(5272) <= inputs(146);
    layer0_outputs(5273) <= not(inputs(245));
    layer0_outputs(5274) <= (inputs(113)) or (inputs(249));
    layer0_outputs(5275) <= (inputs(207)) and not (inputs(132));
    layer0_outputs(5276) <= inputs(247);
    layer0_outputs(5277) <= inputs(87);
    layer0_outputs(5278) <= (inputs(242)) and not (inputs(255));
    layer0_outputs(5279) <= not(inputs(25)) or (inputs(163));
    layer0_outputs(5280) <= '0';
    layer0_outputs(5281) <= not(inputs(71)) or (inputs(34));
    layer0_outputs(5282) <= inputs(6);
    layer0_outputs(5283) <= (inputs(162)) or (inputs(114));
    layer0_outputs(5284) <= '1';
    layer0_outputs(5285) <= '0';
    layer0_outputs(5286) <= not(inputs(210));
    layer0_outputs(5287) <= not(inputs(29)) or (inputs(162));
    layer0_outputs(5288) <= (inputs(106)) and not (inputs(216));
    layer0_outputs(5289) <= (inputs(129)) or (inputs(236));
    layer0_outputs(5290) <= (inputs(254)) and (inputs(116));
    layer0_outputs(5291) <= not(inputs(248));
    layer0_outputs(5292) <= not(inputs(67));
    layer0_outputs(5293) <= inputs(74);
    layer0_outputs(5294) <= inputs(78);
    layer0_outputs(5295) <= not(inputs(237));
    layer0_outputs(5296) <= not(inputs(3)) or (inputs(159));
    layer0_outputs(5297) <= inputs(76);
    layer0_outputs(5298) <= not(inputs(49)) or (inputs(80));
    layer0_outputs(5299) <= (inputs(220)) xor (inputs(114));
    layer0_outputs(5300) <= inputs(135);
    layer0_outputs(5301) <= inputs(138);
    layer0_outputs(5302) <= not(inputs(77));
    layer0_outputs(5303) <= (inputs(43)) or (inputs(37));
    layer0_outputs(5304) <= not(inputs(210));
    layer0_outputs(5305) <= not(inputs(138)) or (inputs(34));
    layer0_outputs(5306) <= not((inputs(45)) xor (inputs(61)));
    layer0_outputs(5307) <= inputs(152);
    layer0_outputs(5308) <= (inputs(23)) or (inputs(203));
    layer0_outputs(5309) <= (inputs(54)) xor (inputs(35));
    layer0_outputs(5310) <= inputs(78);
    layer0_outputs(5311) <= (inputs(93)) or (inputs(95));
    layer0_outputs(5312) <= inputs(61);
    layer0_outputs(5313) <= (inputs(152)) and not (inputs(76));
    layer0_outputs(5314) <= (inputs(27)) and not (inputs(188));
    layer0_outputs(5315) <= not(inputs(43)) or (inputs(239));
    layer0_outputs(5316) <= not(inputs(49)) or (inputs(3));
    layer0_outputs(5317) <= (inputs(46)) and not (inputs(122));
    layer0_outputs(5318) <= not(inputs(72)) or (inputs(159));
    layer0_outputs(5319) <= not(inputs(57)) or (inputs(133));
    layer0_outputs(5320) <= inputs(108);
    layer0_outputs(5321) <= not((inputs(200)) and (inputs(171)));
    layer0_outputs(5322) <= (inputs(210)) or (inputs(221));
    layer0_outputs(5323) <= inputs(223);
    layer0_outputs(5324) <= (inputs(165)) xor (inputs(255));
    layer0_outputs(5325) <= inputs(136);
    layer0_outputs(5326) <= not((inputs(207)) xor (inputs(157)));
    layer0_outputs(5327) <= not(inputs(99));
    layer0_outputs(5328) <= not(inputs(27));
    layer0_outputs(5329) <= (inputs(174)) or (inputs(62));
    layer0_outputs(5330) <= not(inputs(225));
    layer0_outputs(5331) <= inputs(229);
    layer0_outputs(5332) <= not((inputs(12)) and (inputs(129)));
    layer0_outputs(5333) <= inputs(22);
    layer0_outputs(5334) <= not((inputs(203)) xor (inputs(171)));
    layer0_outputs(5335) <= not((inputs(136)) or (inputs(141)));
    layer0_outputs(5336) <= (inputs(46)) or (inputs(104));
    layer0_outputs(5337) <= inputs(161);
    layer0_outputs(5338) <= not((inputs(254)) or (inputs(226)));
    layer0_outputs(5339) <= not(inputs(10)) or (inputs(194));
    layer0_outputs(5340) <= inputs(232);
    layer0_outputs(5341) <= inputs(195);
    layer0_outputs(5342) <= not(inputs(37)) or (inputs(212));
    layer0_outputs(5343) <= not((inputs(103)) or (inputs(168)));
    layer0_outputs(5344) <= not(inputs(124));
    layer0_outputs(5345) <= (inputs(54)) or (inputs(255));
    layer0_outputs(5346) <= not((inputs(37)) or (inputs(96)));
    layer0_outputs(5347) <= not(inputs(230));
    layer0_outputs(5348) <= (inputs(6)) and not (inputs(2));
    layer0_outputs(5349) <= not(inputs(104)) or (inputs(157));
    layer0_outputs(5350) <= (inputs(231)) and not (inputs(151));
    layer0_outputs(5351) <= not((inputs(223)) xor (inputs(177)));
    layer0_outputs(5352) <= inputs(188);
    layer0_outputs(5353) <= not((inputs(111)) xor (inputs(109)));
    layer0_outputs(5354) <= not((inputs(220)) and (inputs(250)));
    layer0_outputs(5355) <= (inputs(195)) xor (inputs(166));
    layer0_outputs(5356) <= (inputs(176)) and not (inputs(252));
    layer0_outputs(5357) <= (inputs(34)) or (inputs(238));
    layer0_outputs(5358) <= inputs(142);
    layer0_outputs(5359) <= not(inputs(228));
    layer0_outputs(5360) <= not(inputs(190));
    layer0_outputs(5361) <= (inputs(221)) xor (inputs(26));
    layer0_outputs(5362) <= '0';
    layer0_outputs(5363) <= not(inputs(64)) or (inputs(68));
    layer0_outputs(5364) <= not(inputs(8));
    layer0_outputs(5365) <= not(inputs(98));
    layer0_outputs(5366) <= not((inputs(229)) or (inputs(6)));
    layer0_outputs(5367) <= (inputs(241)) or (inputs(194));
    layer0_outputs(5368) <= '1';
    layer0_outputs(5369) <= inputs(229);
    layer0_outputs(5370) <= not((inputs(30)) or (inputs(5)));
    layer0_outputs(5371) <= (inputs(141)) or (inputs(222));
    layer0_outputs(5372) <= inputs(233);
    layer0_outputs(5373) <= (inputs(196)) and not (inputs(32));
    layer0_outputs(5374) <= not((inputs(236)) or (inputs(50)));
    layer0_outputs(5375) <= not((inputs(74)) xor (inputs(0)));
    layer0_outputs(5376) <= (inputs(179)) xor (inputs(235));
    layer0_outputs(5377) <= (inputs(170)) xor (inputs(158));
    layer0_outputs(5378) <= not(inputs(178));
    layer0_outputs(5379) <= inputs(249);
    layer0_outputs(5380) <= not((inputs(152)) or (inputs(133)));
    layer0_outputs(5381) <= (inputs(254)) or (inputs(211));
    layer0_outputs(5382) <= (inputs(77)) or (inputs(27));
    layer0_outputs(5383) <= not(inputs(120));
    layer0_outputs(5384) <= not(inputs(180)) or (inputs(16));
    layer0_outputs(5385) <= (inputs(146)) and not (inputs(253));
    layer0_outputs(5386) <= not(inputs(189)) or (inputs(59));
    layer0_outputs(5387) <= (inputs(185)) and not (inputs(235));
    layer0_outputs(5388) <= (inputs(196)) xor (inputs(178));
    layer0_outputs(5389) <= (inputs(107)) and not (inputs(225));
    layer0_outputs(5390) <= not(inputs(246));
    layer0_outputs(5391) <= not(inputs(166)) or (inputs(66));
    layer0_outputs(5392) <= not(inputs(199)) or (inputs(147));
    layer0_outputs(5393) <= (inputs(63)) and not (inputs(242));
    layer0_outputs(5394) <= inputs(152);
    layer0_outputs(5395) <= not(inputs(123)) or (inputs(176));
    layer0_outputs(5396) <= (inputs(115)) and not (inputs(224));
    layer0_outputs(5397) <= not(inputs(238));
    layer0_outputs(5398) <= not(inputs(188));
    layer0_outputs(5399) <= inputs(221);
    layer0_outputs(5400) <= not((inputs(254)) xor (inputs(70)));
    layer0_outputs(5401) <= not(inputs(190)) or (inputs(239));
    layer0_outputs(5402) <= inputs(214);
    layer0_outputs(5403) <= (inputs(189)) or (inputs(171));
    layer0_outputs(5404) <= not((inputs(157)) xor (inputs(192)));
    layer0_outputs(5405) <= not(inputs(194));
    layer0_outputs(5406) <= not((inputs(118)) and (inputs(165)));
    layer0_outputs(5407) <= (inputs(88)) or (inputs(119));
    layer0_outputs(5408) <= not(inputs(20)) or (inputs(86));
    layer0_outputs(5409) <= inputs(91);
    layer0_outputs(5410) <= not(inputs(18)) or (inputs(241));
    layer0_outputs(5411) <= inputs(51);
    layer0_outputs(5412) <= inputs(118);
    layer0_outputs(5413) <= not(inputs(134));
    layer0_outputs(5414) <= inputs(26);
    layer0_outputs(5415) <= (inputs(215)) and not (inputs(251));
    layer0_outputs(5416) <= not((inputs(28)) and (inputs(226)));
    layer0_outputs(5417) <= (inputs(203)) xor (inputs(220));
    layer0_outputs(5418) <= (inputs(106)) and not (inputs(57));
    layer0_outputs(5419) <= not(inputs(112));
    layer0_outputs(5420) <= inputs(153);
    layer0_outputs(5421) <= not(inputs(153)) or (inputs(20));
    layer0_outputs(5422) <= '0';
    layer0_outputs(5423) <= inputs(205);
    layer0_outputs(5424) <= (inputs(25)) and not (inputs(204));
    layer0_outputs(5425) <= not((inputs(84)) or (inputs(202)));
    layer0_outputs(5426) <= not((inputs(200)) or (inputs(206)));
    layer0_outputs(5427) <= not((inputs(40)) or (inputs(33)));
    layer0_outputs(5428) <= inputs(232);
    layer0_outputs(5429) <= not(inputs(106));
    layer0_outputs(5430) <= not(inputs(151)) or (inputs(219));
    layer0_outputs(5431) <= inputs(133);
    layer0_outputs(5432) <= not((inputs(253)) xor (inputs(128)));
    layer0_outputs(5433) <= not((inputs(1)) xor (inputs(223)));
    layer0_outputs(5434) <= not((inputs(242)) or (inputs(33)));
    layer0_outputs(5435) <= inputs(163);
    layer0_outputs(5436) <= not((inputs(237)) xor (inputs(32)));
    layer0_outputs(5437) <= inputs(190);
    layer0_outputs(5438) <= not((inputs(249)) xor (inputs(240)));
    layer0_outputs(5439) <= not((inputs(220)) and (inputs(20)));
    layer0_outputs(5440) <= inputs(122);
    layer0_outputs(5441) <= (inputs(196)) and not (inputs(51));
    layer0_outputs(5442) <= (inputs(63)) or (inputs(124));
    layer0_outputs(5443) <= (inputs(150)) xor (inputs(185));
    layer0_outputs(5444) <= not(inputs(188)) or (inputs(247));
    layer0_outputs(5445) <= not((inputs(218)) xor (inputs(184)));
    layer0_outputs(5446) <= not((inputs(70)) xor (inputs(64)));
    layer0_outputs(5447) <= not((inputs(214)) and (inputs(163)));
    layer0_outputs(5448) <= not(inputs(35)) or (inputs(240));
    layer0_outputs(5449) <= not(inputs(157));
    layer0_outputs(5450) <= not((inputs(74)) or (inputs(44)));
    layer0_outputs(5451) <= (inputs(105)) or (inputs(32));
    layer0_outputs(5452) <= (inputs(138)) and not (inputs(126));
    layer0_outputs(5453) <= (inputs(30)) and not (inputs(253));
    layer0_outputs(5454) <= not(inputs(183));
    layer0_outputs(5455) <= (inputs(68)) xor (inputs(83));
    layer0_outputs(5456) <= (inputs(193)) or (inputs(1));
    layer0_outputs(5457) <= (inputs(81)) and not (inputs(116));
    layer0_outputs(5458) <= inputs(24);
    layer0_outputs(5459) <= (inputs(124)) and (inputs(83));
    layer0_outputs(5460) <= not((inputs(82)) or (inputs(254)));
    layer0_outputs(5461) <= (inputs(245)) and (inputs(175));
    layer0_outputs(5462) <= not((inputs(69)) xor (inputs(18)));
    layer0_outputs(5463) <= (inputs(129)) xor (inputs(86));
    layer0_outputs(5464) <= not(inputs(176)) or (inputs(191));
    layer0_outputs(5465) <= not((inputs(78)) xor (inputs(32)));
    layer0_outputs(5466) <= not(inputs(114)) or (inputs(168));
    layer0_outputs(5467) <= (inputs(58)) and not (inputs(151));
    layer0_outputs(5468) <= '1';
    layer0_outputs(5469) <= not(inputs(217)) or (inputs(240));
    layer0_outputs(5470) <= not(inputs(59));
    layer0_outputs(5471) <= not(inputs(131));
    layer0_outputs(5472) <= (inputs(2)) xor (inputs(172));
    layer0_outputs(5473) <= inputs(108);
    layer0_outputs(5474) <= (inputs(224)) or (inputs(48));
    layer0_outputs(5475) <= (inputs(0)) and not (inputs(2));
    layer0_outputs(5476) <= not(inputs(150)) or (inputs(129));
    layer0_outputs(5477) <= not(inputs(115));
    layer0_outputs(5478) <= (inputs(154)) and not (inputs(51));
    layer0_outputs(5479) <= not(inputs(197)) or (inputs(85));
    layer0_outputs(5480) <= inputs(164);
    layer0_outputs(5481) <= not((inputs(31)) or (inputs(59)));
    layer0_outputs(5482) <= not((inputs(54)) and (inputs(165)));
    layer0_outputs(5483) <= inputs(121);
    layer0_outputs(5484) <= not(inputs(216));
    layer0_outputs(5485) <= not((inputs(202)) xor (inputs(9)));
    layer0_outputs(5486) <= not(inputs(253));
    layer0_outputs(5487) <= inputs(163);
    layer0_outputs(5488) <= inputs(122);
    layer0_outputs(5489) <= (inputs(88)) xor (inputs(212));
    layer0_outputs(5490) <= not((inputs(236)) or (inputs(228)));
    layer0_outputs(5491) <= inputs(27);
    layer0_outputs(5492) <= (inputs(132)) or (inputs(112));
    layer0_outputs(5493) <= (inputs(183)) and not (inputs(199));
    layer0_outputs(5494) <= not(inputs(48)) or (inputs(130));
    layer0_outputs(5495) <= not(inputs(57)) or (inputs(55));
    layer0_outputs(5496) <= (inputs(250)) xor (inputs(220));
    layer0_outputs(5497) <= inputs(135);
    layer0_outputs(5498) <= not((inputs(1)) xor (inputs(186)));
    layer0_outputs(5499) <= not((inputs(253)) xor (inputs(162)));
    layer0_outputs(5500) <= not((inputs(86)) or (inputs(221)));
    layer0_outputs(5501) <= (inputs(212)) or (inputs(112));
    layer0_outputs(5502) <= not((inputs(46)) or (inputs(91)));
    layer0_outputs(5503) <= (inputs(33)) and (inputs(237));
    layer0_outputs(5504) <= '0';
    layer0_outputs(5505) <= not((inputs(211)) and (inputs(94)));
    layer0_outputs(5506) <= not(inputs(174));
    layer0_outputs(5507) <= inputs(194);
    layer0_outputs(5508) <= not(inputs(52));
    layer0_outputs(5509) <= not((inputs(60)) and (inputs(13)));
    layer0_outputs(5510) <= not((inputs(27)) or (inputs(34)));
    layer0_outputs(5511) <= not(inputs(106));
    layer0_outputs(5512) <= inputs(46);
    layer0_outputs(5513) <= not(inputs(130));
    layer0_outputs(5514) <= not(inputs(161)) or (inputs(113));
    layer0_outputs(5515) <= (inputs(194)) or (inputs(214));
    layer0_outputs(5516) <= inputs(82);
    layer0_outputs(5517) <= not(inputs(106));
    layer0_outputs(5518) <= inputs(59);
    layer0_outputs(5519) <= not((inputs(176)) or (inputs(203)));
    layer0_outputs(5520) <= not((inputs(140)) or (inputs(22)));
    layer0_outputs(5521) <= inputs(101);
    layer0_outputs(5522) <= not(inputs(118));
    layer0_outputs(5523) <= (inputs(95)) or (inputs(222));
    layer0_outputs(5524) <= (inputs(173)) and not (inputs(198));
    layer0_outputs(5525) <= not((inputs(88)) or (inputs(190)));
    layer0_outputs(5526) <= (inputs(182)) or (inputs(172));
    layer0_outputs(5527) <= not((inputs(215)) or (inputs(144)));
    layer0_outputs(5528) <= not((inputs(187)) or (inputs(135)));
    layer0_outputs(5529) <= (inputs(96)) or (inputs(184));
    layer0_outputs(5530) <= inputs(106);
    layer0_outputs(5531) <= not((inputs(65)) or (inputs(192)));
    layer0_outputs(5532) <= not(inputs(249));
    layer0_outputs(5533) <= not((inputs(237)) and (inputs(84)));
    layer0_outputs(5534) <= (inputs(24)) or (inputs(35));
    layer0_outputs(5535) <= not((inputs(25)) and (inputs(132)));
    layer0_outputs(5536) <= not((inputs(90)) and (inputs(122)));
    layer0_outputs(5537) <= '1';
    layer0_outputs(5538) <= not(inputs(196));
    layer0_outputs(5539) <= not(inputs(31));
    layer0_outputs(5540) <= not((inputs(36)) xor (inputs(100)));
    layer0_outputs(5541) <= (inputs(110)) or (inputs(127));
    layer0_outputs(5542) <= not((inputs(18)) xor (inputs(5)));
    layer0_outputs(5543) <= not((inputs(2)) xor (inputs(221)));
    layer0_outputs(5544) <= not(inputs(6));
    layer0_outputs(5545) <= not(inputs(164));
    layer0_outputs(5546) <= '1';
    layer0_outputs(5547) <= (inputs(207)) and not (inputs(228));
    layer0_outputs(5548) <= (inputs(77)) and not (inputs(254));
    layer0_outputs(5549) <= (inputs(254)) or (inputs(234));
    layer0_outputs(5550) <= not((inputs(35)) or (inputs(2)));
    layer0_outputs(5551) <= (inputs(38)) and not (inputs(247));
    layer0_outputs(5552) <= (inputs(236)) and not (inputs(56));
    layer0_outputs(5553) <= not(inputs(121)) or (inputs(254));
    layer0_outputs(5554) <= not(inputs(79));
    layer0_outputs(5555) <= inputs(134);
    layer0_outputs(5556) <= inputs(184);
    layer0_outputs(5557) <= inputs(89);
    layer0_outputs(5558) <= (inputs(160)) and (inputs(137));
    layer0_outputs(5559) <= not((inputs(241)) or (inputs(41)));
    layer0_outputs(5560) <= inputs(54);
    layer0_outputs(5561) <= not(inputs(182));
    layer0_outputs(5562) <= not(inputs(197));
    layer0_outputs(5563) <= (inputs(127)) xor (inputs(203));
    layer0_outputs(5564) <= not(inputs(85)) or (inputs(219));
    layer0_outputs(5565) <= (inputs(36)) xor (inputs(118));
    layer0_outputs(5566) <= not(inputs(247)) or (inputs(59));
    layer0_outputs(5567) <= not((inputs(141)) or (inputs(9)));
    layer0_outputs(5568) <= not((inputs(91)) or (inputs(6)));
    layer0_outputs(5569) <= not((inputs(215)) or (inputs(195)));
    layer0_outputs(5570) <= '1';
    layer0_outputs(5571) <= not(inputs(91));
    layer0_outputs(5572) <= not(inputs(142));
    layer0_outputs(5573) <= not((inputs(81)) or (inputs(100)));
    layer0_outputs(5574) <= not(inputs(230));
    layer0_outputs(5575) <= inputs(178);
    layer0_outputs(5576) <= inputs(122);
    layer0_outputs(5577) <= (inputs(24)) xor (inputs(86));
    layer0_outputs(5578) <= '1';
    layer0_outputs(5579) <= (inputs(99)) or (inputs(187));
    layer0_outputs(5580) <= (inputs(39)) and not (inputs(58));
    layer0_outputs(5581) <= inputs(99);
    layer0_outputs(5582) <= inputs(191);
    layer0_outputs(5583) <= not((inputs(252)) xor (inputs(188)));
    layer0_outputs(5584) <= not(inputs(216));
    layer0_outputs(5585) <= not(inputs(102)) or (inputs(56));
    layer0_outputs(5586) <= not(inputs(228)) or (inputs(114));
    layer0_outputs(5587) <= (inputs(34)) and (inputs(73));
    layer0_outputs(5588) <= not(inputs(186));
    layer0_outputs(5589) <= not((inputs(56)) or (inputs(159)));
    layer0_outputs(5590) <= inputs(134);
    layer0_outputs(5591) <= not((inputs(123)) or (inputs(172)));
    layer0_outputs(5592) <= inputs(245);
    layer0_outputs(5593) <= (inputs(19)) xor (inputs(12));
    layer0_outputs(5594) <= not(inputs(107));
    layer0_outputs(5595) <= (inputs(90)) and not (inputs(151));
    layer0_outputs(5596) <= not((inputs(158)) xor (inputs(225)));
    layer0_outputs(5597) <= (inputs(193)) and not (inputs(14));
    layer0_outputs(5598) <= not(inputs(47));
    layer0_outputs(5599) <= not((inputs(174)) or (inputs(224)));
    layer0_outputs(5600) <= inputs(134);
    layer0_outputs(5601) <= (inputs(98)) xor (inputs(101));
    layer0_outputs(5602) <= not((inputs(81)) or (inputs(166)));
    layer0_outputs(5603) <= not((inputs(36)) and (inputs(1)));
    layer0_outputs(5604) <= not((inputs(194)) and (inputs(62)));
    layer0_outputs(5605) <= not(inputs(1)) or (inputs(191));
    layer0_outputs(5606) <= not((inputs(186)) or (inputs(3)));
    layer0_outputs(5607) <= (inputs(180)) and (inputs(168));
    layer0_outputs(5608) <= (inputs(18)) or (inputs(74));
    layer0_outputs(5609) <= (inputs(100)) or (inputs(97));
    layer0_outputs(5610) <= not(inputs(99));
    layer0_outputs(5611) <= (inputs(61)) and (inputs(45));
    layer0_outputs(5612) <= '0';
    layer0_outputs(5613) <= inputs(136);
    layer0_outputs(5614) <= (inputs(178)) and (inputs(41));
    layer0_outputs(5615) <= not(inputs(210));
    layer0_outputs(5616) <= not(inputs(11));
    layer0_outputs(5617) <= inputs(145);
    layer0_outputs(5618) <= (inputs(247)) or (inputs(194));
    layer0_outputs(5619) <= not(inputs(141)) or (inputs(245));
    layer0_outputs(5620) <= '1';
    layer0_outputs(5621) <= not((inputs(152)) or (inputs(182)));
    layer0_outputs(5622) <= not(inputs(191)) or (inputs(238));
    layer0_outputs(5623) <= not((inputs(50)) or (inputs(28)));
    layer0_outputs(5624) <= not((inputs(206)) or (inputs(89)));
    layer0_outputs(5625) <= (inputs(253)) and not (inputs(215));
    layer0_outputs(5626) <= (inputs(98)) or (inputs(172));
    layer0_outputs(5627) <= inputs(174);
    layer0_outputs(5628) <= inputs(40);
    layer0_outputs(5629) <= not((inputs(95)) or (inputs(130)));
    layer0_outputs(5630) <= not((inputs(104)) or (inputs(103)));
    layer0_outputs(5631) <= not(inputs(120)) or (inputs(194));
    layer0_outputs(5632) <= '1';
    layer0_outputs(5633) <= (inputs(242)) or (inputs(38));
    layer0_outputs(5634) <= not(inputs(117));
    layer0_outputs(5635) <= not(inputs(169)) or (inputs(250));
    layer0_outputs(5636) <= not(inputs(101)) or (inputs(4));
    layer0_outputs(5637) <= not(inputs(89));
    layer0_outputs(5638) <= (inputs(244)) and not (inputs(81));
    layer0_outputs(5639) <= not((inputs(252)) or (inputs(24)));
    layer0_outputs(5640) <= (inputs(125)) or (inputs(144));
    layer0_outputs(5641) <= not(inputs(23)) or (inputs(93));
    layer0_outputs(5642) <= (inputs(48)) and not (inputs(126));
    layer0_outputs(5643) <= not(inputs(72)) or (inputs(213));
    layer0_outputs(5644) <= not(inputs(75));
    layer0_outputs(5645) <= inputs(130);
    layer0_outputs(5646) <= (inputs(137)) or (inputs(20));
    layer0_outputs(5647) <= not(inputs(108));
    layer0_outputs(5648) <= inputs(42);
    layer0_outputs(5649) <= inputs(105);
    layer0_outputs(5650) <= (inputs(35)) or (inputs(24));
    layer0_outputs(5651) <= '0';
    layer0_outputs(5652) <= (inputs(182)) xor (inputs(108));
    layer0_outputs(5653) <= not(inputs(160)) or (inputs(200));
    layer0_outputs(5654) <= (inputs(219)) or (inputs(93));
    layer0_outputs(5655) <= not((inputs(120)) and (inputs(23)));
    layer0_outputs(5656) <= (inputs(196)) or (inputs(180));
    layer0_outputs(5657) <= not((inputs(143)) and (inputs(243)));
    layer0_outputs(5658) <= (inputs(234)) or (inputs(104));
    layer0_outputs(5659) <= not(inputs(39));
    layer0_outputs(5660) <= (inputs(37)) and not (inputs(64));
    layer0_outputs(5661) <= not((inputs(17)) xor (inputs(179)));
    layer0_outputs(5662) <= (inputs(123)) and (inputs(3));
    layer0_outputs(5663) <= (inputs(210)) and not (inputs(117));
    layer0_outputs(5664) <= (inputs(123)) and not (inputs(225));
    layer0_outputs(5665) <= (inputs(237)) and (inputs(21));
    layer0_outputs(5666) <= not((inputs(15)) or (inputs(86)));
    layer0_outputs(5667) <= (inputs(156)) and not (inputs(113));
    layer0_outputs(5668) <= not(inputs(136));
    layer0_outputs(5669) <= inputs(166);
    layer0_outputs(5670) <= (inputs(115)) and (inputs(83));
    layer0_outputs(5671) <= inputs(245);
    layer0_outputs(5672) <= (inputs(45)) and not (inputs(90));
    layer0_outputs(5673) <= (inputs(157)) and not (inputs(229));
    layer0_outputs(5674) <= not(inputs(8)) or (inputs(31));
    layer0_outputs(5675) <= not(inputs(254));
    layer0_outputs(5676) <= '0';
    layer0_outputs(5677) <= not(inputs(61)) or (inputs(14));
    layer0_outputs(5678) <= not((inputs(78)) xor (inputs(90)));
    layer0_outputs(5679) <= inputs(86);
    layer0_outputs(5680) <= not((inputs(142)) or (inputs(191)));
    layer0_outputs(5681) <= not((inputs(85)) xor (inputs(205)));
    layer0_outputs(5682) <= inputs(159);
    layer0_outputs(5683) <= not(inputs(101));
    layer0_outputs(5684) <= not((inputs(40)) and (inputs(92)));
    layer0_outputs(5685) <= (inputs(21)) and (inputs(0));
    layer0_outputs(5686) <= (inputs(106)) and (inputs(187));
    layer0_outputs(5687) <= (inputs(63)) or (inputs(39));
    layer0_outputs(5688) <= inputs(174);
    layer0_outputs(5689) <= not((inputs(3)) xor (inputs(62)));
    layer0_outputs(5690) <= not(inputs(37)) or (inputs(220));
    layer0_outputs(5691) <= not(inputs(159)) or (inputs(132));
    layer0_outputs(5692) <= not(inputs(87));
    layer0_outputs(5693) <= (inputs(37)) and not (inputs(239));
    layer0_outputs(5694) <= '1';
    layer0_outputs(5695) <= (inputs(159)) xor (inputs(28));
    layer0_outputs(5696) <= not((inputs(248)) or (inputs(195)));
    layer0_outputs(5697) <= not((inputs(157)) xor (inputs(5)));
    layer0_outputs(5698) <= not((inputs(13)) xor (inputs(232)));
    layer0_outputs(5699) <= not((inputs(51)) or (inputs(23)));
    layer0_outputs(5700) <= not((inputs(115)) or (inputs(148)));
    layer0_outputs(5701) <= (inputs(254)) and not (inputs(35));
    layer0_outputs(5702) <= not(inputs(188));
    layer0_outputs(5703) <= not(inputs(101)) or (inputs(59));
    layer0_outputs(5704) <= '0';
    layer0_outputs(5705) <= (inputs(150)) or (inputs(163));
    layer0_outputs(5706) <= inputs(19);
    layer0_outputs(5707) <= (inputs(122)) xor (inputs(128));
    layer0_outputs(5708) <= inputs(9);
    layer0_outputs(5709) <= not(inputs(143)) or (inputs(30));
    layer0_outputs(5710) <= (inputs(102)) and not (inputs(219));
    layer0_outputs(5711) <= not((inputs(22)) or (inputs(1)));
    layer0_outputs(5712) <= not(inputs(41));
    layer0_outputs(5713) <= not(inputs(103));
    layer0_outputs(5714) <= not(inputs(8));
    layer0_outputs(5715) <= not((inputs(207)) xor (inputs(208)));
    layer0_outputs(5716) <= '1';
    layer0_outputs(5717) <= not((inputs(17)) or (inputs(214)));
    layer0_outputs(5718) <= (inputs(254)) or (inputs(8));
    layer0_outputs(5719) <= not((inputs(98)) or (inputs(56)));
    layer0_outputs(5720) <= (inputs(225)) xor (inputs(132));
    layer0_outputs(5721) <= (inputs(204)) or (inputs(162));
    layer0_outputs(5722) <= not((inputs(80)) or (inputs(203)));
    layer0_outputs(5723) <= (inputs(213)) and not (inputs(75));
    layer0_outputs(5724) <= not(inputs(122));
    layer0_outputs(5725) <= not((inputs(80)) or (inputs(144)));
    layer0_outputs(5726) <= not(inputs(58)) or (inputs(13));
    layer0_outputs(5727) <= (inputs(10)) and not (inputs(218));
    layer0_outputs(5728) <= not(inputs(92));
    layer0_outputs(5729) <= not(inputs(38)) or (inputs(163));
    layer0_outputs(5730) <= not(inputs(100)) or (inputs(55));
    layer0_outputs(5731) <= inputs(103);
    layer0_outputs(5732) <= '0';
    layer0_outputs(5733) <= not((inputs(219)) or (inputs(248)));
    layer0_outputs(5734) <= (inputs(47)) and not (inputs(215));
    layer0_outputs(5735) <= not(inputs(133)) or (inputs(225));
    layer0_outputs(5736) <= inputs(29);
    layer0_outputs(5737) <= not((inputs(119)) or (inputs(133)));
    layer0_outputs(5738) <= not(inputs(218)) or (inputs(118));
    layer0_outputs(5739) <= not(inputs(6)) or (inputs(243));
    layer0_outputs(5740) <= not((inputs(26)) and (inputs(244)));
    layer0_outputs(5741) <= (inputs(212)) and not (inputs(94));
    layer0_outputs(5742) <= (inputs(23)) and not (inputs(238));
    layer0_outputs(5743) <= (inputs(225)) or (inputs(44));
    layer0_outputs(5744) <= '0';
    layer0_outputs(5745) <= (inputs(43)) and (inputs(104));
    layer0_outputs(5746) <= (inputs(37)) and not (inputs(207));
    layer0_outputs(5747) <= (inputs(25)) or (inputs(10));
    layer0_outputs(5748) <= (inputs(211)) and not (inputs(131));
    layer0_outputs(5749) <= (inputs(214)) and (inputs(133));
    layer0_outputs(5750) <= inputs(146);
    layer0_outputs(5751) <= inputs(2);
    layer0_outputs(5752) <= (inputs(234)) and not (inputs(2));
    layer0_outputs(5753) <= not((inputs(36)) and (inputs(71)));
    layer0_outputs(5754) <= not(inputs(228));
    layer0_outputs(5755) <= (inputs(199)) and (inputs(15));
    layer0_outputs(5756) <= inputs(64);
    layer0_outputs(5757) <= not(inputs(247));
    layer0_outputs(5758) <= (inputs(39)) and not (inputs(238));
    layer0_outputs(5759) <= (inputs(32)) and (inputs(80));
    layer0_outputs(5760) <= not((inputs(144)) or (inputs(86)));
    layer0_outputs(5761) <= (inputs(179)) xor (inputs(61));
    layer0_outputs(5762) <= not(inputs(232));
    layer0_outputs(5763) <= not(inputs(44)) or (inputs(119));
    layer0_outputs(5764) <= (inputs(233)) or (inputs(247));
    layer0_outputs(5765) <= not(inputs(120)) or (inputs(41));
    layer0_outputs(5766) <= not(inputs(200));
    layer0_outputs(5767) <= (inputs(28)) xor (inputs(45));
    layer0_outputs(5768) <= not((inputs(46)) or (inputs(55)));
    layer0_outputs(5769) <= not((inputs(104)) xor (inputs(20)));
    layer0_outputs(5770) <= inputs(43);
    layer0_outputs(5771) <= not(inputs(102));
    layer0_outputs(5772) <= not((inputs(156)) xor (inputs(44)));
    layer0_outputs(5773) <= not((inputs(8)) and (inputs(125)));
    layer0_outputs(5774) <= not(inputs(53)) or (inputs(249));
    layer0_outputs(5775) <= not((inputs(210)) xor (inputs(198)));
    layer0_outputs(5776) <= not(inputs(239)) or (inputs(158));
    layer0_outputs(5777) <= (inputs(60)) or (inputs(56));
    layer0_outputs(5778) <= '0';
    layer0_outputs(5779) <= (inputs(242)) and not (inputs(42));
    layer0_outputs(5780) <= not(inputs(221));
    layer0_outputs(5781) <= not((inputs(187)) and (inputs(98)));
    layer0_outputs(5782) <= not(inputs(101)) or (inputs(250));
    layer0_outputs(5783) <= not(inputs(106)) or (inputs(111));
    layer0_outputs(5784) <= (inputs(13)) or (inputs(16));
    layer0_outputs(5785) <= (inputs(249)) and not (inputs(41));
    layer0_outputs(5786) <= not(inputs(23));
    layer0_outputs(5787) <= inputs(0);
    layer0_outputs(5788) <= not(inputs(117));
    layer0_outputs(5789) <= not(inputs(133));
    layer0_outputs(5790) <= not(inputs(67));
    layer0_outputs(5791) <= inputs(150);
    layer0_outputs(5792) <= not((inputs(148)) xor (inputs(117)));
    layer0_outputs(5793) <= not(inputs(240)) or (inputs(199));
    layer0_outputs(5794) <= not(inputs(53)) or (inputs(17));
    layer0_outputs(5795) <= (inputs(120)) xor (inputs(108));
    layer0_outputs(5796) <= not(inputs(89)) or (inputs(162));
    layer0_outputs(5797) <= inputs(193);
    layer0_outputs(5798) <= not((inputs(254)) xor (inputs(247)));
    layer0_outputs(5799) <= not(inputs(74));
    layer0_outputs(5800) <= '1';
    layer0_outputs(5801) <= not((inputs(13)) xor (inputs(82)));
    layer0_outputs(5802) <= '0';
    layer0_outputs(5803) <= (inputs(77)) and not (inputs(165));
    layer0_outputs(5804) <= not(inputs(132));
    layer0_outputs(5805) <= not((inputs(211)) or (inputs(222)));
    layer0_outputs(5806) <= not(inputs(168)) or (inputs(192));
    layer0_outputs(5807) <= not(inputs(40)) or (inputs(113));
    layer0_outputs(5808) <= not((inputs(5)) xor (inputs(136)));
    layer0_outputs(5809) <= (inputs(113)) xor (inputs(240));
    layer0_outputs(5810) <= inputs(138);
    layer0_outputs(5811) <= not(inputs(91)) or (inputs(236));
    layer0_outputs(5812) <= not(inputs(44));
    layer0_outputs(5813) <= '0';
    layer0_outputs(5814) <= (inputs(172)) or (inputs(78));
    layer0_outputs(5815) <= (inputs(105)) xor (inputs(140));
    layer0_outputs(5816) <= (inputs(4)) xor (inputs(122));
    layer0_outputs(5817) <= not((inputs(11)) xor (inputs(174)));
    layer0_outputs(5818) <= not(inputs(229)) or (inputs(89));
    layer0_outputs(5819) <= (inputs(104)) and not (inputs(204));
    layer0_outputs(5820) <= not((inputs(38)) or (inputs(245)));
    layer0_outputs(5821) <= not((inputs(193)) xor (inputs(83)));
    layer0_outputs(5822) <= (inputs(214)) and not (inputs(57));
    layer0_outputs(5823) <= (inputs(115)) or (inputs(149));
    layer0_outputs(5824) <= not(inputs(97));
    layer0_outputs(5825) <= not((inputs(255)) and (inputs(223)));
    layer0_outputs(5826) <= not(inputs(217));
    layer0_outputs(5827) <= not(inputs(73)) or (inputs(179));
    layer0_outputs(5828) <= not((inputs(149)) and (inputs(244)));
    layer0_outputs(5829) <= not(inputs(26));
    layer0_outputs(5830) <= (inputs(156)) xor (inputs(218));
    layer0_outputs(5831) <= not((inputs(131)) and (inputs(131)));
    layer0_outputs(5832) <= not(inputs(27)) or (inputs(218));
    layer0_outputs(5833) <= not(inputs(75));
    layer0_outputs(5834) <= not((inputs(238)) or (inputs(219)));
    layer0_outputs(5835) <= not(inputs(205));
    layer0_outputs(5836) <= (inputs(88)) and not (inputs(206));
    layer0_outputs(5837) <= (inputs(130)) and not (inputs(29));
    layer0_outputs(5838) <= not(inputs(54));
    layer0_outputs(5839) <= inputs(174);
    layer0_outputs(5840) <= inputs(56);
    layer0_outputs(5841) <= not((inputs(131)) or (inputs(135)));
    layer0_outputs(5842) <= inputs(93);
    layer0_outputs(5843) <= not(inputs(36));
    layer0_outputs(5844) <= not(inputs(24));
    layer0_outputs(5845) <= (inputs(62)) and (inputs(106));
    layer0_outputs(5846) <= inputs(76);
    layer0_outputs(5847) <= (inputs(39)) or (inputs(45));
    layer0_outputs(5848) <= (inputs(214)) or (inputs(196));
    layer0_outputs(5849) <= (inputs(241)) or (inputs(61));
    layer0_outputs(5850) <= not(inputs(169));
    layer0_outputs(5851) <= not((inputs(35)) or (inputs(15)));
    layer0_outputs(5852) <= not((inputs(250)) and (inputs(200)));
    layer0_outputs(5853) <= not(inputs(115));
    layer0_outputs(5854) <= not(inputs(154)) or (inputs(194));
    layer0_outputs(5855) <= inputs(193);
    layer0_outputs(5856) <= (inputs(123)) and (inputs(194));
    layer0_outputs(5857) <= inputs(9);
    layer0_outputs(5858) <= (inputs(225)) and not (inputs(93));
    layer0_outputs(5859) <= not((inputs(191)) xor (inputs(193)));
    layer0_outputs(5860) <= not(inputs(39));
    layer0_outputs(5861) <= not(inputs(153)) or (inputs(39));
    layer0_outputs(5862) <= not(inputs(232)) or (inputs(46));
    layer0_outputs(5863) <= not(inputs(180));
    layer0_outputs(5864) <= not(inputs(145));
    layer0_outputs(5865) <= inputs(185);
    layer0_outputs(5866) <= not(inputs(215)) or (inputs(41));
    layer0_outputs(5867) <= not(inputs(67)) or (inputs(13));
    layer0_outputs(5868) <= not((inputs(255)) or (inputs(14)));
    layer0_outputs(5869) <= (inputs(38)) or (inputs(115));
    layer0_outputs(5870) <= not((inputs(244)) and (inputs(248)));
    layer0_outputs(5871) <= inputs(186);
    layer0_outputs(5872) <= not((inputs(202)) or (inputs(224)));
    layer0_outputs(5873) <= not(inputs(127));
    layer0_outputs(5874) <= not((inputs(191)) xor (inputs(49)));
    layer0_outputs(5875) <= inputs(64);
    layer0_outputs(5876) <= not((inputs(59)) or (inputs(4)));
    layer0_outputs(5877) <= '1';
    layer0_outputs(5878) <= not((inputs(252)) or (inputs(250)));
    layer0_outputs(5879) <= not(inputs(16)) or (inputs(59));
    layer0_outputs(5880) <= (inputs(2)) and not (inputs(65));
    layer0_outputs(5881) <= not(inputs(97)) or (inputs(41));
    layer0_outputs(5882) <= (inputs(23)) xor (inputs(60));
    layer0_outputs(5883) <= not(inputs(206)) or (inputs(213));
    layer0_outputs(5884) <= not((inputs(201)) or (inputs(67)));
    layer0_outputs(5885) <= '0';
    layer0_outputs(5886) <= not((inputs(135)) or (inputs(35)));
    layer0_outputs(5887) <= not(inputs(132)) or (inputs(65));
    layer0_outputs(5888) <= (inputs(229)) and not (inputs(110));
    layer0_outputs(5889) <= (inputs(60)) or (inputs(165));
    layer0_outputs(5890) <= not((inputs(194)) or (inputs(191)));
    layer0_outputs(5891) <= '0';
    layer0_outputs(5892) <= '0';
    layer0_outputs(5893) <= not(inputs(25));
    layer0_outputs(5894) <= (inputs(69)) or (inputs(239));
    layer0_outputs(5895) <= '0';
    layer0_outputs(5896) <= not(inputs(212)) or (inputs(192));
    layer0_outputs(5897) <= not((inputs(146)) xor (inputs(85)));
    layer0_outputs(5898) <= (inputs(134)) and not (inputs(20));
    layer0_outputs(5899) <= not((inputs(24)) and (inputs(27)));
    layer0_outputs(5900) <= not(inputs(54));
    layer0_outputs(5901) <= '0';
    layer0_outputs(5902) <= (inputs(248)) and not (inputs(191));
    layer0_outputs(5903) <= not(inputs(122));
    layer0_outputs(5904) <= inputs(70);
    layer0_outputs(5905) <= '0';
    layer0_outputs(5906) <= (inputs(16)) or (inputs(110));
    layer0_outputs(5907) <= (inputs(37)) or (inputs(5));
    layer0_outputs(5908) <= not(inputs(233));
    layer0_outputs(5909) <= (inputs(243)) or (inputs(70));
    layer0_outputs(5910) <= inputs(247);
    layer0_outputs(5911) <= '1';
    layer0_outputs(5912) <= not(inputs(201));
    layer0_outputs(5913) <= (inputs(171)) or (inputs(102));
    layer0_outputs(5914) <= inputs(193);
    layer0_outputs(5915) <= inputs(83);
    layer0_outputs(5916) <= not(inputs(180)) or (inputs(80));
    layer0_outputs(5917) <= not(inputs(211));
    layer0_outputs(5918) <= inputs(180);
    layer0_outputs(5919) <= (inputs(39)) and (inputs(78));
    layer0_outputs(5920) <= (inputs(9)) and not (inputs(72));
    layer0_outputs(5921) <= not(inputs(112));
    layer0_outputs(5922) <= inputs(103);
    layer0_outputs(5923) <= not(inputs(204)) or (inputs(225));
    layer0_outputs(5924) <= inputs(45);
    layer0_outputs(5925) <= not(inputs(198)) or (inputs(47));
    layer0_outputs(5926) <= not((inputs(210)) and (inputs(117)));
    layer0_outputs(5927) <= not((inputs(157)) or (inputs(243)));
    layer0_outputs(5928) <= not(inputs(160)) or (inputs(186));
    layer0_outputs(5929) <= '1';
    layer0_outputs(5930) <= not(inputs(246)) or (inputs(213));
    layer0_outputs(5931) <= not((inputs(194)) or (inputs(127)));
    layer0_outputs(5932) <= not(inputs(127));
    layer0_outputs(5933) <= (inputs(98)) xor (inputs(121));
    layer0_outputs(5934) <= not(inputs(246)) or (inputs(241));
    layer0_outputs(5935) <= (inputs(193)) and not (inputs(146));
    layer0_outputs(5936) <= not(inputs(55)) or (inputs(204));
    layer0_outputs(5937) <= (inputs(134)) and not (inputs(191));
    layer0_outputs(5938) <= inputs(90);
    layer0_outputs(5939) <= inputs(58);
    layer0_outputs(5940) <= inputs(217);
    layer0_outputs(5941) <= not(inputs(192)) or (inputs(6));
    layer0_outputs(5942) <= inputs(9);
    layer0_outputs(5943) <= inputs(65);
    layer0_outputs(5944) <= (inputs(165)) or (inputs(66));
    layer0_outputs(5945) <= inputs(203);
    layer0_outputs(5946) <= '1';
    layer0_outputs(5947) <= inputs(56);
    layer0_outputs(5948) <= inputs(104);
    layer0_outputs(5949) <= not(inputs(162)) or (inputs(76));
    layer0_outputs(5950) <= not(inputs(110));
    layer0_outputs(5951) <= (inputs(210)) and not (inputs(120));
    layer0_outputs(5952) <= (inputs(36)) xor (inputs(67));
    layer0_outputs(5953) <= '1';
    layer0_outputs(5954) <= not(inputs(54));
    layer0_outputs(5955) <= not((inputs(96)) and (inputs(32)));
    layer0_outputs(5956) <= inputs(203);
    layer0_outputs(5957) <= not(inputs(180)) or (inputs(13));
    layer0_outputs(5958) <= inputs(153);
    layer0_outputs(5959) <= not(inputs(92));
    layer0_outputs(5960) <= not((inputs(86)) xor (inputs(66)));
    layer0_outputs(5961) <= not(inputs(57)) or (inputs(97));
    layer0_outputs(5962) <= (inputs(176)) or (inputs(95));
    layer0_outputs(5963) <= (inputs(169)) or (inputs(233));
    layer0_outputs(5964) <= (inputs(159)) and not (inputs(94));
    layer0_outputs(5965) <= inputs(87);
    layer0_outputs(5966) <= (inputs(82)) or (inputs(191));
    layer0_outputs(5967) <= '0';
    layer0_outputs(5968) <= (inputs(177)) or (inputs(70));
    layer0_outputs(5969) <= inputs(154);
    layer0_outputs(5970) <= '0';
    layer0_outputs(5971) <= (inputs(196)) and (inputs(8));
    layer0_outputs(5972) <= inputs(59);
    layer0_outputs(5973) <= not(inputs(133)) or (inputs(39));
    layer0_outputs(5974) <= (inputs(232)) or (inputs(96));
    layer0_outputs(5975) <= not((inputs(206)) or (inputs(33)));
    layer0_outputs(5976) <= (inputs(97)) or (inputs(53));
    layer0_outputs(5977) <= not((inputs(161)) or (inputs(144)));
    layer0_outputs(5978) <= inputs(139);
    layer0_outputs(5979) <= not((inputs(124)) xor (inputs(155)));
    layer0_outputs(5980) <= not(inputs(54));
    layer0_outputs(5981) <= not(inputs(220)) or (inputs(200));
    layer0_outputs(5982) <= not(inputs(84));
    layer0_outputs(5983) <= not(inputs(49));
    layer0_outputs(5984) <= not(inputs(68));
    layer0_outputs(5985) <= (inputs(100)) and not (inputs(72));
    layer0_outputs(5986) <= (inputs(174)) or (inputs(42));
    layer0_outputs(5987) <= not(inputs(220)) or (inputs(15));
    layer0_outputs(5988) <= (inputs(115)) and (inputs(195));
    layer0_outputs(5989) <= inputs(104);
    layer0_outputs(5990) <= not(inputs(218)) or (inputs(174));
    layer0_outputs(5991) <= not(inputs(187));
    layer0_outputs(5992) <= not(inputs(99));
    layer0_outputs(5993) <= inputs(165);
    layer0_outputs(5994) <= inputs(160);
    layer0_outputs(5995) <= (inputs(251)) xor (inputs(243));
    layer0_outputs(5996) <= not(inputs(30));
    layer0_outputs(5997) <= not(inputs(31)) or (inputs(99));
    layer0_outputs(5998) <= not(inputs(227));
    layer0_outputs(5999) <= not((inputs(133)) xor (inputs(176)));
    layer0_outputs(6000) <= not(inputs(39));
    layer0_outputs(6001) <= (inputs(117)) and not (inputs(3));
    layer0_outputs(6002) <= not(inputs(105));
    layer0_outputs(6003) <= (inputs(27)) and (inputs(208));
    layer0_outputs(6004) <= not((inputs(114)) xor (inputs(63)));
    layer0_outputs(6005) <= not(inputs(199));
    layer0_outputs(6006) <= not((inputs(203)) xor (inputs(170)));
    layer0_outputs(6007) <= not(inputs(59));
    layer0_outputs(6008) <= (inputs(94)) and not (inputs(149));
    layer0_outputs(6009) <= not((inputs(58)) or (inputs(142)));
    layer0_outputs(6010) <= '1';
    layer0_outputs(6011) <= inputs(111);
    layer0_outputs(6012) <= not((inputs(185)) xor (inputs(1)));
    layer0_outputs(6013) <= inputs(206);
    layer0_outputs(6014) <= not((inputs(23)) or (inputs(94)));
    layer0_outputs(6015) <= inputs(64);
    layer0_outputs(6016) <= inputs(52);
    layer0_outputs(6017) <= not(inputs(69));
    layer0_outputs(6018) <= (inputs(200)) and not (inputs(97));
    layer0_outputs(6019) <= inputs(90);
    layer0_outputs(6020) <= '0';
    layer0_outputs(6021) <= not(inputs(44)) or (inputs(221));
    layer0_outputs(6022) <= not(inputs(227));
    layer0_outputs(6023) <= inputs(26);
    layer0_outputs(6024) <= inputs(129);
    layer0_outputs(6025) <= not(inputs(211)) or (inputs(253));
    layer0_outputs(6026) <= not(inputs(185));
    layer0_outputs(6027) <= (inputs(65)) and not (inputs(124));
    layer0_outputs(6028) <= not(inputs(201));
    layer0_outputs(6029) <= '1';
    layer0_outputs(6030) <= '0';
    layer0_outputs(6031) <= not(inputs(186));
    layer0_outputs(6032) <= inputs(181);
    layer0_outputs(6033) <= not(inputs(5)) or (inputs(146));
    layer0_outputs(6034) <= inputs(0);
    layer0_outputs(6035) <= inputs(236);
    layer0_outputs(6036) <= not(inputs(101));
    layer0_outputs(6037) <= (inputs(233)) and not (inputs(90));
    layer0_outputs(6038) <= (inputs(56)) and not (inputs(152));
    layer0_outputs(6039) <= not(inputs(187)) or (inputs(97));
    layer0_outputs(6040) <= not((inputs(226)) xor (inputs(65)));
    layer0_outputs(6041) <= (inputs(7)) or (inputs(244));
    layer0_outputs(6042) <= not(inputs(238));
    layer0_outputs(6043) <= (inputs(229)) and (inputs(147));
    layer0_outputs(6044) <= (inputs(191)) or (inputs(187));
    layer0_outputs(6045) <= (inputs(117)) or (inputs(45));
    layer0_outputs(6046) <= not(inputs(183)) or (inputs(96));
    layer0_outputs(6047) <= inputs(164);
    layer0_outputs(6048) <= not(inputs(181)) or (inputs(58));
    layer0_outputs(6049) <= (inputs(82)) or (inputs(54));
    layer0_outputs(6050) <= not((inputs(104)) xor (inputs(21)));
    layer0_outputs(6051) <= inputs(57);
    layer0_outputs(6052) <= not(inputs(110));
    layer0_outputs(6053) <= not(inputs(216));
    layer0_outputs(6054) <= (inputs(7)) and not (inputs(247));
    layer0_outputs(6055) <= not((inputs(206)) and (inputs(74)));
    layer0_outputs(6056) <= not(inputs(148));
    layer0_outputs(6057) <= not(inputs(212)) or (inputs(46));
    layer0_outputs(6058) <= inputs(27);
    layer0_outputs(6059) <= not(inputs(248));
    layer0_outputs(6060) <= '1';
    layer0_outputs(6061) <= (inputs(241)) and not (inputs(128));
    layer0_outputs(6062) <= (inputs(157)) or (inputs(185));
    layer0_outputs(6063) <= not(inputs(233)) or (inputs(181));
    layer0_outputs(6064) <= (inputs(53)) or (inputs(209));
    layer0_outputs(6065) <= not(inputs(227));
    layer0_outputs(6066) <= '0';
    layer0_outputs(6067) <= not(inputs(228)) or (inputs(152));
    layer0_outputs(6068) <= '0';
    layer0_outputs(6069) <= not((inputs(176)) xor (inputs(23)));
    layer0_outputs(6070) <= inputs(24);
    layer0_outputs(6071) <= inputs(203);
    layer0_outputs(6072) <= (inputs(37)) and not (inputs(71));
    layer0_outputs(6073) <= (inputs(245)) and (inputs(87));
    layer0_outputs(6074) <= (inputs(220)) and not (inputs(58));
    layer0_outputs(6075) <= not(inputs(152));
    layer0_outputs(6076) <= not((inputs(102)) or (inputs(39)));
    layer0_outputs(6077) <= not(inputs(234));
    layer0_outputs(6078) <= (inputs(249)) xor (inputs(185));
    layer0_outputs(6079) <= not(inputs(229));
    layer0_outputs(6080) <= not(inputs(197));
    layer0_outputs(6081) <= not(inputs(2));
    layer0_outputs(6082) <= not((inputs(28)) and (inputs(78)));
    layer0_outputs(6083) <= not(inputs(185)) or (inputs(98));
    layer0_outputs(6084) <= inputs(22);
    layer0_outputs(6085) <= not(inputs(44));
    layer0_outputs(6086) <= not((inputs(87)) and (inputs(23)));
    layer0_outputs(6087) <= not(inputs(20));
    layer0_outputs(6088) <= not(inputs(213)) or (inputs(157));
    layer0_outputs(6089) <= not(inputs(0)) or (inputs(81));
    layer0_outputs(6090) <= not(inputs(30));
    layer0_outputs(6091) <= not(inputs(53)) or (inputs(0));
    layer0_outputs(6092) <= not((inputs(171)) xor (inputs(205)));
    layer0_outputs(6093) <= not((inputs(34)) xor (inputs(108)));
    layer0_outputs(6094) <= inputs(142);
    layer0_outputs(6095) <= '0';
    layer0_outputs(6096) <= not(inputs(18)) or (inputs(113));
    layer0_outputs(6097) <= not(inputs(243)) or (inputs(131));
    layer0_outputs(6098) <= not((inputs(197)) or (inputs(158)));
    layer0_outputs(6099) <= '0';
    layer0_outputs(6100) <= (inputs(88)) or (inputs(187));
    layer0_outputs(6101) <= not(inputs(83));
    layer0_outputs(6102) <= inputs(176);
    layer0_outputs(6103) <= not(inputs(255)) or (inputs(150));
    layer0_outputs(6104) <= not(inputs(166));
    layer0_outputs(6105) <= not(inputs(74));
    layer0_outputs(6106) <= not(inputs(24)) or (inputs(143));
    layer0_outputs(6107) <= inputs(70);
    layer0_outputs(6108) <= not(inputs(9)) or (inputs(14));
    layer0_outputs(6109) <= (inputs(57)) and (inputs(46));
    layer0_outputs(6110) <= not(inputs(49));
    layer0_outputs(6111) <= not((inputs(63)) or (inputs(10)));
    layer0_outputs(6112) <= inputs(181);
    layer0_outputs(6113) <= (inputs(152)) and not (inputs(126));
    layer0_outputs(6114) <= not(inputs(168));
    layer0_outputs(6115) <= (inputs(62)) and not (inputs(129));
    layer0_outputs(6116) <= (inputs(114)) xor (inputs(86));
    layer0_outputs(6117) <= not(inputs(220));
    layer0_outputs(6118) <= not((inputs(227)) xor (inputs(197)));
    layer0_outputs(6119) <= not(inputs(156)) or (inputs(6));
    layer0_outputs(6120) <= inputs(148);
    layer0_outputs(6121) <= not(inputs(231)) or (inputs(121));
    layer0_outputs(6122) <= (inputs(151)) or (inputs(238));
    layer0_outputs(6123) <= not(inputs(117));
    layer0_outputs(6124) <= (inputs(248)) or (inputs(132));
    layer0_outputs(6125) <= not(inputs(136));
    layer0_outputs(6126) <= inputs(49);
    layer0_outputs(6127) <= inputs(137);
    layer0_outputs(6128) <= not((inputs(194)) or (inputs(193)));
    layer0_outputs(6129) <= (inputs(99)) or (inputs(213));
    layer0_outputs(6130) <= not(inputs(67));
    layer0_outputs(6131) <= not(inputs(198));
    layer0_outputs(6132) <= inputs(23);
    layer0_outputs(6133) <= (inputs(31)) or (inputs(59));
    layer0_outputs(6134) <= (inputs(164)) and not (inputs(1));
    layer0_outputs(6135) <= not((inputs(162)) or (inputs(219)));
    layer0_outputs(6136) <= not(inputs(94));
    layer0_outputs(6137) <= not((inputs(106)) or (inputs(144)));
    layer0_outputs(6138) <= not(inputs(115)) or (inputs(16));
    layer0_outputs(6139) <= not((inputs(244)) xor (inputs(165)));
    layer0_outputs(6140) <= not(inputs(124)) or (inputs(71));
    layer0_outputs(6141) <= (inputs(213)) and (inputs(125));
    layer0_outputs(6142) <= (inputs(197)) and (inputs(96));
    layer0_outputs(6143) <= not((inputs(63)) or (inputs(25)));
    layer0_outputs(6144) <= not((inputs(133)) or (inputs(133)));
    layer0_outputs(6145) <= (inputs(159)) or (inputs(199));
    layer0_outputs(6146) <= inputs(47);
    layer0_outputs(6147) <= not(inputs(210)) or (inputs(96));
    layer0_outputs(6148) <= not(inputs(213));
    layer0_outputs(6149) <= not(inputs(28)) or (inputs(118));
    layer0_outputs(6150) <= (inputs(106)) xor (inputs(102));
    layer0_outputs(6151) <= not((inputs(150)) or (inputs(185)));
    layer0_outputs(6152) <= not(inputs(107));
    layer0_outputs(6153) <= not((inputs(69)) or (inputs(246)));
    layer0_outputs(6154) <= inputs(79);
    layer0_outputs(6155) <= not(inputs(70)) or (inputs(19));
    layer0_outputs(6156) <= not(inputs(138));
    layer0_outputs(6157) <= not(inputs(230));
    layer0_outputs(6158) <= (inputs(235)) xor (inputs(186));
    layer0_outputs(6159) <= not(inputs(56));
    layer0_outputs(6160) <= not(inputs(156));
    layer0_outputs(6161) <= (inputs(105)) xor (inputs(93));
    layer0_outputs(6162) <= not((inputs(188)) and (inputs(218)));
    layer0_outputs(6163) <= (inputs(160)) xor (inputs(147));
    layer0_outputs(6164) <= not((inputs(216)) and (inputs(43)));
    layer0_outputs(6165) <= not((inputs(181)) xor (inputs(228)));
    layer0_outputs(6166) <= not(inputs(136));
    layer0_outputs(6167) <= not((inputs(249)) xor (inputs(217)));
    layer0_outputs(6168) <= not(inputs(214)) or (inputs(105));
    layer0_outputs(6169) <= (inputs(105)) or (inputs(183));
    layer0_outputs(6170) <= inputs(36);
    layer0_outputs(6171) <= not((inputs(27)) or (inputs(143)));
    layer0_outputs(6172) <= (inputs(52)) or (inputs(68));
    layer0_outputs(6173) <= not((inputs(173)) xor (inputs(170)));
    layer0_outputs(6174) <= not((inputs(122)) and (inputs(79)));
    layer0_outputs(6175) <= not((inputs(136)) or (inputs(142)));
    layer0_outputs(6176) <= inputs(197);
    layer0_outputs(6177) <= (inputs(168)) and not (inputs(61));
    layer0_outputs(6178) <= (inputs(90)) or (inputs(180));
    layer0_outputs(6179) <= not(inputs(108)) or (inputs(229));
    layer0_outputs(6180) <= (inputs(176)) or (inputs(235));
    layer0_outputs(6181) <= not(inputs(115));
    layer0_outputs(6182) <= not((inputs(242)) xor (inputs(144)));
    layer0_outputs(6183) <= (inputs(132)) and (inputs(147));
    layer0_outputs(6184) <= not(inputs(49)) or (inputs(253));
    layer0_outputs(6185) <= not(inputs(88));
    layer0_outputs(6186) <= (inputs(140)) and not (inputs(209));
    layer0_outputs(6187) <= not((inputs(249)) and (inputs(199)));
    layer0_outputs(6188) <= inputs(152);
    layer0_outputs(6189) <= inputs(54);
    layer0_outputs(6190) <= not(inputs(217));
    layer0_outputs(6191) <= (inputs(235)) xor (inputs(191));
    layer0_outputs(6192) <= (inputs(20)) and (inputs(183));
    layer0_outputs(6193) <= not(inputs(96));
    layer0_outputs(6194) <= not(inputs(110)) or (inputs(95));
    layer0_outputs(6195) <= not(inputs(54));
    layer0_outputs(6196) <= not(inputs(77)) or (inputs(253));
    layer0_outputs(6197) <= '0';
    layer0_outputs(6198) <= not(inputs(228)) or (inputs(182));
    layer0_outputs(6199) <= (inputs(52)) and not (inputs(252));
    layer0_outputs(6200) <= inputs(92);
    layer0_outputs(6201) <= not((inputs(216)) or (inputs(191)));
    layer0_outputs(6202) <= (inputs(236)) or (inputs(4));
    layer0_outputs(6203) <= (inputs(119)) and not (inputs(24));
    layer0_outputs(6204) <= not((inputs(48)) or (inputs(207)));
    layer0_outputs(6205) <= not((inputs(167)) or (inputs(83)));
    layer0_outputs(6206) <= not(inputs(134));
    layer0_outputs(6207) <= (inputs(162)) and not (inputs(240));
    layer0_outputs(6208) <= not(inputs(197)) or (inputs(34));
    layer0_outputs(6209) <= not(inputs(47)) or (inputs(170));
    layer0_outputs(6210) <= not(inputs(100)) or (inputs(207));
    layer0_outputs(6211) <= inputs(3);
    layer0_outputs(6212) <= (inputs(191)) or (inputs(134));
    layer0_outputs(6213) <= not(inputs(101));
    layer0_outputs(6214) <= not(inputs(196));
    layer0_outputs(6215) <= (inputs(170)) xor (inputs(85));
    layer0_outputs(6216) <= inputs(117);
    layer0_outputs(6217) <= not(inputs(44));
    layer0_outputs(6218) <= inputs(68);
    layer0_outputs(6219) <= inputs(121);
    layer0_outputs(6220) <= (inputs(55)) and (inputs(126));
    layer0_outputs(6221) <= not(inputs(104));
    layer0_outputs(6222) <= not((inputs(161)) or (inputs(212)));
    layer0_outputs(6223) <= (inputs(149)) and not (inputs(60));
    layer0_outputs(6224) <= (inputs(49)) and not (inputs(189));
    layer0_outputs(6225) <= (inputs(172)) and not (inputs(168));
    layer0_outputs(6226) <= (inputs(64)) and (inputs(119));
    layer0_outputs(6227) <= not((inputs(239)) or (inputs(137)));
    layer0_outputs(6228) <= not(inputs(92));
    layer0_outputs(6229) <= (inputs(92)) xor (inputs(51));
    layer0_outputs(6230) <= not(inputs(17));
    layer0_outputs(6231) <= inputs(163);
    layer0_outputs(6232) <= inputs(64);
    layer0_outputs(6233) <= not(inputs(197)) or (inputs(156));
    layer0_outputs(6234) <= inputs(41);
    layer0_outputs(6235) <= inputs(57);
    layer0_outputs(6236) <= (inputs(108)) xor (inputs(3));
    layer0_outputs(6237) <= not(inputs(119)) or (inputs(0));
    layer0_outputs(6238) <= (inputs(125)) and (inputs(146));
    layer0_outputs(6239) <= inputs(104);
    layer0_outputs(6240) <= (inputs(40)) and not (inputs(102));
    layer0_outputs(6241) <= not((inputs(120)) or (inputs(118)));
    layer0_outputs(6242) <= not(inputs(108));
    layer0_outputs(6243) <= (inputs(229)) or (inputs(139));
    layer0_outputs(6244) <= not((inputs(120)) xor (inputs(217)));
    layer0_outputs(6245) <= not(inputs(52));
    layer0_outputs(6246) <= not(inputs(25)) or (inputs(215));
    layer0_outputs(6247) <= not((inputs(150)) or (inputs(14)));
    layer0_outputs(6248) <= not(inputs(19)) or (inputs(192));
    layer0_outputs(6249) <= inputs(241);
    layer0_outputs(6250) <= (inputs(186)) and not (inputs(86));
    layer0_outputs(6251) <= inputs(114);
    layer0_outputs(6252) <= not((inputs(96)) or (inputs(230)));
    layer0_outputs(6253) <= not((inputs(220)) or (inputs(239)));
    layer0_outputs(6254) <= not(inputs(179));
    layer0_outputs(6255) <= (inputs(220)) or (inputs(169));
    layer0_outputs(6256) <= (inputs(74)) and not (inputs(223));
    layer0_outputs(6257) <= not(inputs(162));
    layer0_outputs(6258) <= not(inputs(170));
    layer0_outputs(6259) <= not((inputs(9)) and (inputs(69)));
    layer0_outputs(6260) <= (inputs(178)) and not (inputs(142));
    layer0_outputs(6261) <= '1';
    layer0_outputs(6262) <= (inputs(125)) or (inputs(99));
    layer0_outputs(6263) <= not(inputs(138));
    layer0_outputs(6264) <= inputs(249);
    layer0_outputs(6265) <= not(inputs(127));
    layer0_outputs(6266) <= inputs(52);
    layer0_outputs(6267) <= not(inputs(110)) or (inputs(199));
    layer0_outputs(6268) <= (inputs(100)) and not (inputs(189));
    layer0_outputs(6269) <= inputs(177);
    layer0_outputs(6270) <= (inputs(5)) or (inputs(183));
    layer0_outputs(6271) <= '0';
    layer0_outputs(6272) <= not((inputs(144)) or (inputs(220)));
    layer0_outputs(6273) <= not(inputs(29));
    layer0_outputs(6274) <= not(inputs(78)) or (inputs(47));
    layer0_outputs(6275) <= not(inputs(213));
    layer0_outputs(6276) <= (inputs(141)) or (inputs(45));
    layer0_outputs(6277) <= (inputs(73)) xor (inputs(141));
    layer0_outputs(6278) <= not((inputs(125)) and (inputs(240)));
    layer0_outputs(6279) <= (inputs(158)) xor (inputs(131));
    layer0_outputs(6280) <= not(inputs(61)) or (inputs(175));
    layer0_outputs(6281) <= not((inputs(204)) xor (inputs(225)));
    layer0_outputs(6282) <= not((inputs(68)) or (inputs(226)));
    layer0_outputs(6283) <= (inputs(44)) and not (inputs(163));
    layer0_outputs(6284) <= (inputs(155)) and not (inputs(167));
    layer0_outputs(6285) <= (inputs(209)) xor (inputs(176));
    layer0_outputs(6286) <= inputs(10);
    layer0_outputs(6287) <= not(inputs(132)) or (inputs(26));
    layer0_outputs(6288) <= not(inputs(116));
    layer0_outputs(6289) <= not((inputs(17)) xor (inputs(89)));
    layer0_outputs(6290) <= inputs(107);
    layer0_outputs(6291) <= (inputs(119)) or (inputs(242));
    layer0_outputs(6292) <= inputs(167);
    layer0_outputs(6293) <= not(inputs(80));
    layer0_outputs(6294) <= (inputs(253)) or (inputs(243));
    layer0_outputs(6295) <= (inputs(30)) and not (inputs(156));
    layer0_outputs(6296) <= not((inputs(132)) or (inputs(226)));
    layer0_outputs(6297) <= not((inputs(231)) or (inputs(180)));
    layer0_outputs(6298) <= not(inputs(13)) or (inputs(55));
    layer0_outputs(6299) <= not(inputs(119));
    layer0_outputs(6300) <= not((inputs(114)) or (inputs(114)));
    layer0_outputs(6301) <= not(inputs(181));
    layer0_outputs(6302) <= not(inputs(134)) or (inputs(116));
    layer0_outputs(6303) <= (inputs(181)) and not (inputs(241));
    layer0_outputs(6304) <= not(inputs(109));
    layer0_outputs(6305) <= not(inputs(165)) or (inputs(134));
    layer0_outputs(6306) <= inputs(66);
    layer0_outputs(6307) <= not((inputs(36)) or (inputs(23)));
    layer0_outputs(6308) <= inputs(102);
    layer0_outputs(6309) <= (inputs(17)) or (inputs(225));
    layer0_outputs(6310) <= not(inputs(22)) or (inputs(98));
    layer0_outputs(6311) <= not((inputs(221)) or (inputs(112)));
    layer0_outputs(6312) <= (inputs(169)) and not (inputs(198));
    layer0_outputs(6313) <= '0';
    layer0_outputs(6314) <= (inputs(80)) xor (inputs(253));
    layer0_outputs(6315) <= (inputs(30)) and not (inputs(212));
    layer0_outputs(6316) <= not(inputs(181));
    layer0_outputs(6317) <= not((inputs(60)) or (inputs(68)));
    layer0_outputs(6318) <= inputs(191);
    layer0_outputs(6319) <= (inputs(205)) or (inputs(147));
    layer0_outputs(6320) <= inputs(154);
    layer0_outputs(6321) <= not((inputs(133)) xor (inputs(162)));
    layer0_outputs(6322) <= (inputs(21)) and not (inputs(130));
    layer0_outputs(6323) <= '1';
    layer0_outputs(6324) <= (inputs(234)) or (inputs(242));
    layer0_outputs(6325) <= not((inputs(106)) or (inputs(206)));
    layer0_outputs(6326) <= (inputs(68)) and not (inputs(208));
    layer0_outputs(6327) <= not(inputs(4));
    layer0_outputs(6328) <= (inputs(154)) or (inputs(189));
    layer0_outputs(6329) <= inputs(238);
    layer0_outputs(6330) <= not(inputs(23));
    layer0_outputs(6331) <= inputs(189);
    layer0_outputs(6332) <= not(inputs(245)) or (inputs(124));
    layer0_outputs(6333) <= inputs(95);
    layer0_outputs(6334) <= not(inputs(136));
    layer0_outputs(6335) <= not((inputs(34)) or (inputs(46)));
    layer0_outputs(6336) <= (inputs(250)) or (inputs(253));
    layer0_outputs(6337) <= not((inputs(221)) xor (inputs(141)));
    layer0_outputs(6338) <= (inputs(88)) xor (inputs(171));
    layer0_outputs(6339) <= (inputs(213)) xor (inputs(66));
    layer0_outputs(6340) <= not((inputs(15)) or (inputs(233)));
    layer0_outputs(6341) <= inputs(157);
    layer0_outputs(6342) <= not((inputs(150)) or (inputs(133)));
    layer0_outputs(6343) <= not(inputs(207));
    layer0_outputs(6344) <= not((inputs(222)) or (inputs(208)));
    layer0_outputs(6345) <= not(inputs(115)) or (inputs(124));
    layer0_outputs(6346) <= not((inputs(81)) xor (inputs(109)));
    layer0_outputs(6347) <= (inputs(170)) or (inputs(143));
    layer0_outputs(6348) <= inputs(179);
    layer0_outputs(6349) <= not((inputs(104)) or (inputs(152)));
    layer0_outputs(6350) <= inputs(246);
    layer0_outputs(6351) <= (inputs(34)) or (inputs(19));
    layer0_outputs(6352) <= (inputs(229)) and not (inputs(72));
    layer0_outputs(6353) <= (inputs(227)) and not (inputs(208));
    layer0_outputs(6354) <= (inputs(61)) and not (inputs(224));
    layer0_outputs(6355) <= not(inputs(131));
    layer0_outputs(6356) <= not(inputs(172));
    layer0_outputs(6357) <= inputs(254);
    layer0_outputs(6358) <= not(inputs(207));
    layer0_outputs(6359) <= not((inputs(223)) or (inputs(219)));
    layer0_outputs(6360) <= '0';
    layer0_outputs(6361) <= not((inputs(170)) or (inputs(7)));
    layer0_outputs(6362) <= (inputs(210)) and (inputs(70));
    layer0_outputs(6363) <= (inputs(251)) xor (inputs(207));
    layer0_outputs(6364) <= inputs(108);
    layer0_outputs(6365) <= (inputs(115)) and not (inputs(224));
    layer0_outputs(6366) <= inputs(151);
    layer0_outputs(6367) <= inputs(15);
    layer0_outputs(6368) <= inputs(131);
    layer0_outputs(6369) <= not((inputs(255)) xor (inputs(98)));
    layer0_outputs(6370) <= not((inputs(129)) and (inputs(230)));
    layer0_outputs(6371) <= not(inputs(182));
    layer0_outputs(6372) <= not(inputs(230));
    layer0_outputs(6373) <= inputs(122);
    layer0_outputs(6374) <= inputs(68);
    layer0_outputs(6375) <= not(inputs(233)) or (inputs(241));
    layer0_outputs(6376) <= not(inputs(240));
    layer0_outputs(6377) <= (inputs(253)) xor (inputs(167));
    layer0_outputs(6378) <= not(inputs(149));
    layer0_outputs(6379) <= (inputs(65)) xor (inputs(87));
    layer0_outputs(6380) <= inputs(135);
    layer0_outputs(6381) <= not((inputs(221)) or (inputs(119)));
    layer0_outputs(6382) <= (inputs(15)) xor (inputs(234));
    layer0_outputs(6383) <= not((inputs(114)) xor (inputs(135)));
    layer0_outputs(6384) <= not((inputs(182)) or (inputs(205)));
    layer0_outputs(6385) <= (inputs(163)) xor (inputs(186));
    layer0_outputs(6386) <= not((inputs(69)) or (inputs(150)));
    layer0_outputs(6387) <= inputs(206);
    layer0_outputs(6388) <= inputs(62);
    layer0_outputs(6389) <= not((inputs(139)) or (inputs(158)));
    layer0_outputs(6390) <= not((inputs(246)) or (inputs(115)));
    layer0_outputs(6391) <= (inputs(69)) and not (inputs(109));
    layer0_outputs(6392) <= not((inputs(70)) xor (inputs(68)));
    layer0_outputs(6393) <= not(inputs(35));
    layer0_outputs(6394) <= not((inputs(240)) and (inputs(48)));
    layer0_outputs(6395) <= inputs(113);
    layer0_outputs(6396) <= not(inputs(34)) or (inputs(129));
    layer0_outputs(6397) <= (inputs(62)) or (inputs(189));
    layer0_outputs(6398) <= (inputs(140)) and not (inputs(211));
    layer0_outputs(6399) <= inputs(75);
    layer0_outputs(6400) <= '1';
    layer0_outputs(6401) <= inputs(53);
    layer0_outputs(6402) <= not((inputs(45)) or (inputs(22)));
    layer0_outputs(6403) <= not((inputs(106)) or (inputs(92)));
    layer0_outputs(6404) <= (inputs(70)) and not (inputs(149));
    layer0_outputs(6405) <= not(inputs(7)) or (inputs(218));
    layer0_outputs(6406) <= (inputs(169)) xor (inputs(189));
    layer0_outputs(6407) <= (inputs(9)) or (inputs(42));
    layer0_outputs(6408) <= not((inputs(250)) and (inputs(170)));
    layer0_outputs(6409) <= not((inputs(51)) or (inputs(52)));
    layer0_outputs(6410) <= not((inputs(149)) xor (inputs(222)));
    layer0_outputs(6411) <= not((inputs(97)) xor (inputs(188)));
    layer0_outputs(6412) <= (inputs(17)) xor (inputs(48));
    layer0_outputs(6413) <= not(inputs(142));
    layer0_outputs(6414) <= (inputs(163)) or (inputs(165));
    layer0_outputs(6415) <= not((inputs(114)) or (inputs(234)));
    layer0_outputs(6416) <= inputs(89);
    layer0_outputs(6417) <= not(inputs(21)) or (inputs(150));
    layer0_outputs(6418) <= not(inputs(114));
    layer0_outputs(6419) <= (inputs(163)) xor (inputs(190));
    layer0_outputs(6420) <= not((inputs(78)) or (inputs(50)));
    layer0_outputs(6421) <= (inputs(237)) xor (inputs(190));
    layer0_outputs(6422) <= not((inputs(31)) xor (inputs(183)));
    layer0_outputs(6423) <= (inputs(134)) and not (inputs(55));
    layer0_outputs(6424) <= not(inputs(151)) or (inputs(185));
    layer0_outputs(6425) <= not(inputs(165));
    layer0_outputs(6426) <= '1';
    layer0_outputs(6427) <= not((inputs(195)) xor (inputs(30)));
    layer0_outputs(6428) <= inputs(153);
    layer0_outputs(6429) <= not((inputs(17)) xor (inputs(222)));
    layer0_outputs(6430) <= '1';
    layer0_outputs(6431) <= not(inputs(215));
    layer0_outputs(6432) <= not(inputs(208)) or (inputs(17));
    layer0_outputs(6433) <= not(inputs(182));
    layer0_outputs(6434) <= (inputs(5)) or (inputs(207));
    layer0_outputs(6435) <= (inputs(33)) or (inputs(98));
    layer0_outputs(6436) <= (inputs(216)) or (inputs(80));
    layer0_outputs(6437) <= (inputs(34)) xor (inputs(238));
    layer0_outputs(6438) <= (inputs(236)) or (inputs(114));
    layer0_outputs(6439) <= not((inputs(9)) or (inputs(144)));
    layer0_outputs(6440) <= not(inputs(39));
    layer0_outputs(6441) <= not((inputs(218)) and (inputs(148)));
    layer0_outputs(6442) <= not(inputs(2)) or (inputs(42));
    layer0_outputs(6443) <= '0';
    layer0_outputs(6444) <= not((inputs(112)) xor (inputs(36)));
    layer0_outputs(6445) <= inputs(106);
    layer0_outputs(6446) <= (inputs(75)) xor (inputs(147));
    layer0_outputs(6447) <= inputs(171);
    layer0_outputs(6448) <= not(inputs(174));
    layer0_outputs(6449) <= not(inputs(8)) or (inputs(138));
    layer0_outputs(6450) <= not(inputs(160));
    layer0_outputs(6451) <= (inputs(187)) and not (inputs(86));
    layer0_outputs(6452) <= (inputs(3)) and not (inputs(114));
    layer0_outputs(6453) <= (inputs(194)) and not (inputs(0));
    layer0_outputs(6454) <= (inputs(10)) or (inputs(147));
    layer0_outputs(6455) <= (inputs(193)) or (inputs(179));
    layer0_outputs(6456) <= not((inputs(213)) or (inputs(218)));
    layer0_outputs(6457) <= not((inputs(151)) or (inputs(252)));
    layer0_outputs(6458) <= not(inputs(39));
    layer0_outputs(6459) <= (inputs(121)) and (inputs(131));
    layer0_outputs(6460) <= inputs(160);
    layer0_outputs(6461) <= not((inputs(32)) or (inputs(172)));
    layer0_outputs(6462) <= inputs(234);
    layer0_outputs(6463) <= not(inputs(101));
    layer0_outputs(6464) <= inputs(255);
    layer0_outputs(6465) <= not((inputs(149)) and (inputs(75)));
    layer0_outputs(6466) <= '0';
    layer0_outputs(6467) <= not(inputs(212));
    layer0_outputs(6468) <= (inputs(74)) and (inputs(111));
    layer0_outputs(6469) <= (inputs(93)) xor (inputs(20));
    layer0_outputs(6470) <= '1';
    layer0_outputs(6471) <= inputs(161);
    layer0_outputs(6472) <= '1';
    layer0_outputs(6473) <= inputs(126);
    layer0_outputs(6474) <= inputs(209);
    layer0_outputs(6475) <= inputs(29);
    layer0_outputs(6476) <= not(inputs(99));
    layer0_outputs(6477) <= not((inputs(150)) or (inputs(79)));
    layer0_outputs(6478) <= not(inputs(112));
    layer0_outputs(6479) <= not((inputs(51)) or (inputs(216)));
    layer0_outputs(6480) <= (inputs(210)) and not (inputs(40));
    layer0_outputs(6481) <= '0';
    layer0_outputs(6482) <= not(inputs(198)) or (inputs(42));
    layer0_outputs(6483) <= (inputs(24)) xor (inputs(26));
    layer0_outputs(6484) <= (inputs(89)) and not (inputs(203));
    layer0_outputs(6485) <= inputs(84);
    layer0_outputs(6486) <= not((inputs(212)) and (inputs(155)));
    layer0_outputs(6487) <= '1';
    layer0_outputs(6488) <= inputs(237);
    layer0_outputs(6489) <= not((inputs(33)) and (inputs(13)));
    layer0_outputs(6490) <= not(inputs(24)) or (inputs(72));
    layer0_outputs(6491) <= '1';
    layer0_outputs(6492) <= (inputs(127)) or (inputs(160));
    layer0_outputs(6493) <= (inputs(137)) xor (inputs(0));
    layer0_outputs(6494) <= (inputs(233)) or (inputs(87));
    layer0_outputs(6495) <= (inputs(62)) and not (inputs(249));
    layer0_outputs(6496) <= (inputs(119)) or (inputs(89));
    layer0_outputs(6497) <= not(inputs(88));
    layer0_outputs(6498) <= not((inputs(100)) or (inputs(10)));
    layer0_outputs(6499) <= not(inputs(87)) or (inputs(194));
    layer0_outputs(6500) <= '1';
    layer0_outputs(6501) <= inputs(37);
    layer0_outputs(6502) <= (inputs(25)) or (inputs(102));
    layer0_outputs(6503) <= (inputs(185)) or (inputs(53));
    layer0_outputs(6504) <= not((inputs(164)) and (inputs(234)));
    layer0_outputs(6505) <= (inputs(201)) and not (inputs(226));
    layer0_outputs(6506) <= not((inputs(192)) xor (inputs(192)));
    layer0_outputs(6507) <= (inputs(30)) and (inputs(242));
    layer0_outputs(6508) <= not(inputs(184));
    layer0_outputs(6509) <= (inputs(154)) or (inputs(214));
    layer0_outputs(6510) <= (inputs(114)) and not (inputs(14));
    layer0_outputs(6511) <= not(inputs(172)) or (inputs(90));
    layer0_outputs(6512) <= not((inputs(90)) xor (inputs(119)));
    layer0_outputs(6513) <= not(inputs(190));
    layer0_outputs(6514) <= not(inputs(220)) or (inputs(126));
    layer0_outputs(6515) <= not(inputs(227));
    layer0_outputs(6516) <= not(inputs(89)) or (inputs(140));
    layer0_outputs(6517) <= not(inputs(102));
    layer0_outputs(6518) <= not((inputs(189)) or (inputs(142)));
    layer0_outputs(6519) <= not(inputs(220));
    layer0_outputs(6520) <= (inputs(157)) xor (inputs(48));
    layer0_outputs(6521) <= not(inputs(219));
    layer0_outputs(6522) <= not((inputs(197)) or (inputs(163)));
    layer0_outputs(6523) <= (inputs(186)) xor (inputs(3));
    layer0_outputs(6524) <= not((inputs(193)) or (inputs(156)));
    layer0_outputs(6525) <= (inputs(119)) and (inputs(69));
    layer0_outputs(6526) <= not((inputs(102)) and (inputs(96)));
    layer0_outputs(6527) <= not(inputs(19)) or (inputs(244));
    layer0_outputs(6528) <= not(inputs(153));
    layer0_outputs(6529) <= (inputs(79)) xor (inputs(236));
    layer0_outputs(6530) <= not(inputs(47));
    layer0_outputs(6531) <= (inputs(15)) and (inputs(125));
    layer0_outputs(6532) <= '1';
    layer0_outputs(6533) <= not((inputs(102)) xor (inputs(128)));
    layer0_outputs(6534) <= not(inputs(195));
    layer0_outputs(6535) <= '1';
    layer0_outputs(6536) <= not(inputs(77));
    layer0_outputs(6537) <= (inputs(67)) and not (inputs(24));
    layer0_outputs(6538) <= not(inputs(230));
    layer0_outputs(6539) <= (inputs(64)) or (inputs(178));
    layer0_outputs(6540) <= inputs(127);
    layer0_outputs(6541) <= (inputs(239)) or (inputs(64));
    layer0_outputs(6542) <= not(inputs(125));
    layer0_outputs(6543) <= inputs(231);
    layer0_outputs(6544) <= not(inputs(19));
    layer0_outputs(6545) <= (inputs(30)) and not (inputs(143));
    layer0_outputs(6546) <= not(inputs(116)) or (inputs(31));
    layer0_outputs(6547) <= not((inputs(128)) or (inputs(113)));
    layer0_outputs(6548) <= not((inputs(70)) or (inputs(112)));
    layer0_outputs(6549) <= not(inputs(143));
    layer0_outputs(6550) <= inputs(237);
    layer0_outputs(6551) <= (inputs(92)) and not (inputs(114));
    layer0_outputs(6552) <= not((inputs(95)) or (inputs(63)));
    layer0_outputs(6553) <= not((inputs(36)) or (inputs(165)));
    layer0_outputs(6554) <= (inputs(157)) or (inputs(6));
    layer0_outputs(6555) <= not((inputs(69)) or (inputs(246)));
    layer0_outputs(6556) <= not(inputs(151)) or (inputs(64));
    layer0_outputs(6557) <= inputs(112);
    layer0_outputs(6558) <= inputs(104);
    layer0_outputs(6559) <= not((inputs(221)) or (inputs(215)));
    layer0_outputs(6560) <= (inputs(247)) or (inputs(145));
    layer0_outputs(6561) <= (inputs(167)) and not (inputs(248));
    layer0_outputs(6562) <= not(inputs(231));
    layer0_outputs(6563) <= not(inputs(126)) or (inputs(198));
    layer0_outputs(6564) <= not(inputs(33));
    layer0_outputs(6565) <= inputs(124);
    layer0_outputs(6566) <= inputs(55);
    layer0_outputs(6567) <= (inputs(124)) and not (inputs(240));
    layer0_outputs(6568) <= not(inputs(166)) or (inputs(78));
    layer0_outputs(6569) <= not(inputs(117));
    layer0_outputs(6570) <= '0';
    layer0_outputs(6571) <= not((inputs(22)) or (inputs(64)));
    layer0_outputs(6572) <= not((inputs(78)) or (inputs(238)));
    layer0_outputs(6573) <= (inputs(194)) or (inputs(201));
    layer0_outputs(6574) <= not(inputs(67)) or (inputs(142));
    layer0_outputs(6575) <= not((inputs(248)) or (inputs(65)));
    layer0_outputs(6576) <= not(inputs(141)) or (inputs(3));
    layer0_outputs(6577) <= not(inputs(106));
    layer0_outputs(6578) <= inputs(8);
    layer0_outputs(6579) <= inputs(78);
    layer0_outputs(6580) <= not(inputs(247)) or (inputs(63));
    layer0_outputs(6581) <= not((inputs(5)) xor (inputs(155)));
    layer0_outputs(6582) <= inputs(81);
    layer0_outputs(6583) <= not(inputs(214));
    layer0_outputs(6584) <= inputs(25);
    layer0_outputs(6585) <= (inputs(139)) and (inputs(48));
    layer0_outputs(6586) <= not(inputs(104));
    layer0_outputs(6587) <= not(inputs(193));
    layer0_outputs(6588) <= (inputs(248)) xor (inputs(170));
    layer0_outputs(6589) <= not(inputs(200));
    layer0_outputs(6590) <= not((inputs(210)) and (inputs(231)));
    layer0_outputs(6591) <= not((inputs(226)) or (inputs(14)));
    layer0_outputs(6592) <= not((inputs(192)) xor (inputs(94)));
    layer0_outputs(6593) <= not(inputs(114));
    layer0_outputs(6594) <= not((inputs(113)) xor (inputs(24)));
    layer0_outputs(6595) <= not(inputs(162)) or (inputs(29));
    layer0_outputs(6596) <= inputs(130);
    layer0_outputs(6597) <= inputs(104);
    layer0_outputs(6598) <= (inputs(201)) or (inputs(231));
    layer0_outputs(6599) <= not(inputs(61));
    layer0_outputs(6600) <= not((inputs(139)) or (inputs(154)));
    layer0_outputs(6601) <= inputs(213);
    layer0_outputs(6602) <= inputs(61);
    layer0_outputs(6603) <= not(inputs(57)) or (inputs(171));
    layer0_outputs(6604) <= inputs(40);
    layer0_outputs(6605) <= inputs(91);
    layer0_outputs(6606) <= not(inputs(123));
    layer0_outputs(6607) <= inputs(228);
    layer0_outputs(6608) <= inputs(143);
    layer0_outputs(6609) <= not((inputs(227)) xor (inputs(254)));
    layer0_outputs(6610) <= inputs(42);
    layer0_outputs(6611) <= (inputs(21)) and not (inputs(144));
    layer0_outputs(6612) <= not(inputs(14));
    layer0_outputs(6613) <= (inputs(24)) or (inputs(48));
    layer0_outputs(6614) <= not((inputs(241)) and (inputs(199)));
    layer0_outputs(6615) <= not((inputs(175)) or (inputs(48)));
    layer0_outputs(6616) <= inputs(66);
    layer0_outputs(6617) <= not(inputs(21)) or (inputs(162));
    layer0_outputs(6618) <= not((inputs(161)) or (inputs(205)));
    layer0_outputs(6619) <= not(inputs(176));
    layer0_outputs(6620) <= (inputs(119)) and not (inputs(237));
    layer0_outputs(6621) <= (inputs(157)) or (inputs(157));
    layer0_outputs(6622) <= not(inputs(226));
    layer0_outputs(6623) <= not(inputs(146));
    layer0_outputs(6624) <= (inputs(5)) or (inputs(106));
    layer0_outputs(6625) <= (inputs(48)) xor (inputs(14));
    layer0_outputs(6626) <= not((inputs(221)) or (inputs(32)));
    layer0_outputs(6627) <= not(inputs(214)) or (inputs(81));
    layer0_outputs(6628) <= inputs(206);
    layer0_outputs(6629) <= (inputs(238)) or (inputs(219));
    layer0_outputs(6630) <= not(inputs(165));
    layer0_outputs(6631) <= not((inputs(44)) or (inputs(50)));
    layer0_outputs(6632) <= not((inputs(146)) or (inputs(44)));
    layer0_outputs(6633) <= '0';
    layer0_outputs(6634) <= inputs(216);
    layer0_outputs(6635) <= (inputs(152)) and not (inputs(22));
    layer0_outputs(6636) <= inputs(55);
    layer0_outputs(6637) <= (inputs(130)) or (inputs(181));
    layer0_outputs(6638) <= (inputs(206)) or (inputs(246));
    layer0_outputs(6639) <= inputs(98);
    layer0_outputs(6640) <= (inputs(97)) or (inputs(230));
    layer0_outputs(6641) <= (inputs(113)) or (inputs(126));
    layer0_outputs(6642) <= inputs(135);
    layer0_outputs(6643) <= '1';
    layer0_outputs(6644) <= not((inputs(190)) or (inputs(14)));
    layer0_outputs(6645) <= inputs(98);
    layer0_outputs(6646) <= (inputs(122)) and not (inputs(49));
    layer0_outputs(6647) <= not(inputs(25));
    layer0_outputs(6648) <= inputs(180);
    layer0_outputs(6649) <= not(inputs(58));
    layer0_outputs(6650) <= inputs(91);
    layer0_outputs(6651) <= (inputs(82)) xor (inputs(72));
    layer0_outputs(6652) <= not(inputs(82));
    layer0_outputs(6653) <= (inputs(198)) and (inputs(96));
    layer0_outputs(6654) <= not((inputs(97)) or (inputs(251)));
    layer0_outputs(6655) <= inputs(247);
    layer0_outputs(6656) <= not(inputs(106));
    layer0_outputs(6657) <= (inputs(34)) and not (inputs(239));
    layer0_outputs(6658) <= not(inputs(162));
    layer0_outputs(6659) <= inputs(82);
    layer0_outputs(6660) <= inputs(153);
    layer0_outputs(6661) <= (inputs(60)) or (inputs(27));
    layer0_outputs(6662) <= (inputs(130)) xor (inputs(101));
    layer0_outputs(6663) <= (inputs(55)) xor (inputs(8));
    layer0_outputs(6664) <= '0';
    layer0_outputs(6665) <= (inputs(135)) or (inputs(243));
    layer0_outputs(6666) <= not(inputs(114));
    layer0_outputs(6667) <= not((inputs(99)) xor (inputs(21)));
    layer0_outputs(6668) <= not(inputs(167)) or (inputs(63));
    layer0_outputs(6669) <= inputs(157);
    layer0_outputs(6670) <= inputs(66);
    layer0_outputs(6671) <= (inputs(239)) or (inputs(180));
    layer0_outputs(6672) <= inputs(249);
    layer0_outputs(6673) <= not(inputs(233));
    layer0_outputs(6674) <= not(inputs(161));
    layer0_outputs(6675) <= not((inputs(165)) or (inputs(181)));
    layer0_outputs(6676) <= (inputs(52)) and not (inputs(27));
    layer0_outputs(6677) <= inputs(104);
    layer0_outputs(6678) <= not(inputs(116));
    layer0_outputs(6679) <= (inputs(108)) and not (inputs(207));
    layer0_outputs(6680) <= not(inputs(39));
    layer0_outputs(6681) <= (inputs(6)) and not (inputs(27));
    layer0_outputs(6682) <= not(inputs(137));
    layer0_outputs(6683) <= not(inputs(188)) or (inputs(122));
    layer0_outputs(6684) <= (inputs(137)) and not (inputs(101));
    layer0_outputs(6685) <= not(inputs(87));
    layer0_outputs(6686) <= not((inputs(141)) and (inputs(137)));
    layer0_outputs(6687) <= inputs(126);
    layer0_outputs(6688) <= not((inputs(10)) or (inputs(106)));
    layer0_outputs(6689) <= not((inputs(71)) xor (inputs(226)));
    layer0_outputs(6690) <= (inputs(110)) or (inputs(12));
    layer0_outputs(6691) <= inputs(16);
    layer0_outputs(6692) <= inputs(130);
    layer0_outputs(6693) <= not(inputs(232)) or (inputs(33));
    layer0_outputs(6694) <= not((inputs(19)) xor (inputs(26)));
    layer0_outputs(6695) <= not(inputs(123)) or (inputs(142));
    layer0_outputs(6696) <= (inputs(135)) and not (inputs(17));
    layer0_outputs(6697) <= inputs(86);
    layer0_outputs(6698) <= inputs(24);
    layer0_outputs(6699) <= inputs(210);
    layer0_outputs(6700) <= not((inputs(55)) or (inputs(116)));
    layer0_outputs(6701) <= not(inputs(75));
    layer0_outputs(6702) <= not((inputs(120)) and (inputs(170)));
    layer0_outputs(6703) <= inputs(164);
    layer0_outputs(6704) <= (inputs(246)) and not (inputs(255));
    layer0_outputs(6705) <= '1';
    layer0_outputs(6706) <= not(inputs(36));
    layer0_outputs(6707) <= (inputs(103)) and not (inputs(16));
    layer0_outputs(6708) <= (inputs(154)) and not (inputs(108));
    layer0_outputs(6709) <= '0';
    layer0_outputs(6710) <= (inputs(80)) or (inputs(60));
    layer0_outputs(6711) <= not(inputs(134)) or (inputs(232));
    layer0_outputs(6712) <= not((inputs(183)) and (inputs(219)));
    layer0_outputs(6713) <= not((inputs(30)) or (inputs(14)));
    layer0_outputs(6714) <= inputs(175);
    layer0_outputs(6715) <= (inputs(192)) and not (inputs(236));
    layer0_outputs(6716) <= inputs(167);
    layer0_outputs(6717) <= (inputs(147)) xor (inputs(100));
    layer0_outputs(6718) <= not((inputs(6)) or (inputs(80)));
    layer0_outputs(6719) <= (inputs(220)) or (inputs(227));
    layer0_outputs(6720) <= (inputs(173)) and (inputs(152));
    layer0_outputs(6721) <= not((inputs(20)) and (inputs(20)));
    layer0_outputs(6722) <= (inputs(121)) and (inputs(56));
    layer0_outputs(6723) <= (inputs(20)) or (inputs(1));
    layer0_outputs(6724) <= (inputs(169)) and not (inputs(53));
    layer0_outputs(6725) <= (inputs(210)) or (inputs(82));
    layer0_outputs(6726) <= not(inputs(120)) or (inputs(204));
    layer0_outputs(6727) <= not((inputs(189)) or (inputs(82)));
    layer0_outputs(6728) <= inputs(119);
    layer0_outputs(6729) <= inputs(219);
    layer0_outputs(6730) <= (inputs(136)) xor (inputs(98));
    layer0_outputs(6731) <= not((inputs(45)) xor (inputs(51)));
    layer0_outputs(6732) <= (inputs(4)) or (inputs(199));
    layer0_outputs(6733) <= (inputs(208)) or (inputs(78));
    layer0_outputs(6734) <= not((inputs(80)) or (inputs(115)));
    layer0_outputs(6735) <= not(inputs(201));
    layer0_outputs(6736) <= inputs(36);
    layer0_outputs(6737) <= not((inputs(252)) or (inputs(106)));
    layer0_outputs(6738) <= not((inputs(70)) or (inputs(178)));
    layer0_outputs(6739) <= (inputs(213)) and (inputs(39));
    layer0_outputs(6740) <= not((inputs(202)) or (inputs(41)));
    layer0_outputs(6741) <= not(inputs(240));
    layer0_outputs(6742) <= not((inputs(98)) or (inputs(128)));
    layer0_outputs(6743) <= not((inputs(120)) and (inputs(60)));
    layer0_outputs(6744) <= not(inputs(43));
    layer0_outputs(6745) <= not(inputs(233));
    layer0_outputs(6746) <= not(inputs(79)) or (inputs(200));
    layer0_outputs(6747) <= '1';
    layer0_outputs(6748) <= not((inputs(109)) or (inputs(82)));
    layer0_outputs(6749) <= (inputs(221)) and not (inputs(30));
    layer0_outputs(6750) <= (inputs(94)) and not (inputs(1));
    layer0_outputs(6751) <= not((inputs(197)) and (inputs(81)));
    layer0_outputs(6752) <= (inputs(62)) and not (inputs(248));
    layer0_outputs(6753) <= not((inputs(57)) and (inputs(39)));
    layer0_outputs(6754) <= not(inputs(76));
    layer0_outputs(6755) <= not((inputs(156)) or (inputs(43)));
    layer0_outputs(6756) <= not((inputs(82)) or (inputs(49)));
    layer0_outputs(6757) <= not((inputs(245)) or (inputs(34)));
    layer0_outputs(6758) <= (inputs(178)) and not (inputs(113));
    layer0_outputs(6759) <= '1';
    layer0_outputs(6760) <= not((inputs(192)) xor (inputs(254)));
    layer0_outputs(6761) <= not((inputs(30)) or (inputs(209)));
    layer0_outputs(6762) <= inputs(139);
    layer0_outputs(6763) <= not(inputs(99));
    layer0_outputs(6764) <= (inputs(126)) or (inputs(14));
    layer0_outputs(6765) <= (inputs(57)) or (inputs(162));
    layer0_outputs(6766) <= inputs(241);
    layer0_outputs(6767) <= inputs(186);
    layer0_outputs(6768) <= not(inputs(49));
    layer0_outputs(6769) <= (inputs(93)) and (inputs(157));
    layer0_outputs(6770) <= (inputs(224)) xor (inputs(152));
    layer0_outputs(6771) <= inputs(191);
    layer0_outputs(6772) <= (inputs(53)) and not (inputs(213));
    layer0_outputs(6773) <= inputs(192);
    layer0_outputs(6774) <= not(inputs(125));
    layer0_outputs(6775) <= not(inputs(83)) or (inputs(208));
    layer0_outputs(6776) <= (inputs(77)) and (inputs(69));
    layer0_outputs(6777) <= not(inputs(155)) or (inputs(19));
    layer0_outputs(6778) <= inputs(222);
    layer0_outputs(6779) <= not(inputs(187));
    layer0_outputs(6780) <= not(inputs(73));
    layer0_outputs(6781) <= (inputs(248)) and (inputs(243));
    layer0_outputs(6782) <= not((inputs(1)) xor (inputs(61)));
    layer0_outputs(6783) <= not((inputs(251)) and (inputs(93)));
    layer0_outputs(6784) <= inputs(21);
    layer0_outputs(6785) <= (inputs(250)) and not (inputs(85));
    layer0_outputs(6786) <= (inputs(120)) xor (inputs(107));
    layer0_outputs(6787) <= not((inputs(220)) xor (inputs(190)));
    layer0_outputs(6788) <= (inputs(202)) and not (inputs(81));
    layer0_outputs(6789) <= not(inputs(229));
    layer0_outputs(6790) <= inputs(137);
    layer0_outputs(6791) <= not(inputs(231));
    layer0_outputs(6792) <= not((inputs(201)) or (inputs(11)));
    layer0_outputs(6793) <= (inputs(106)) and not (inputs(181));
    layer0_outputs(6794) <= not((inputs(112)) xor (inputs(129)));
    layer0_outputs(6795) <= not(inputs(36)) or (inputs(160));
    layer0_outputs(6796) <= not(inputs(7)) or (inputs(23));
    layer0_outputs(6797) <= inputs(254);
    layer0_outputs(6798) <= (inputs(84)) or (inputs(155));
    layer0_outputs(6799) <= not(inputs(161));
    layer0_outputs(6800) <= (inputs(57)) and not (inputs(162));
    layer0_outputs(6801) <= (inputs(82)) or (inputs(116));
    layer0_outputs(6802) <= '0';
    layer0_outputs(6803) <= not(inputs(203)) or (inputs(30));
    layer0_outputs(6804) <= not(inputs(89));
    layer0_outputs(6805) <= not(inputs(188));
    layer0_outputs(6806) <= not(inputs(159));
    layer0_outputs(6807) <= not(inputs(162)) or (inputs(248));
    layer0_outputs(6808) <= not(inputs(1));
    layer0_outputs(6809) <= not(inputs(203)) or (inputs(70));
    layer0_outputs(6810) <= inputs(151);
    layer0_outputs(6811) <= not((inputs(254)) xor (inputs(147)));
    layer0_outputs(6812) <= not(inputs(114));
    layer0_outputs(6813) <= not(inputs(98));
    layer0_outputs(6814) <= not(inputs(67));
    layer0_outputs(6815) <= not(inputs(92));
    layer0_outputs(6816) <= not((inputs(145)) or (inputs(84)));
    layer0_outputs(6817) <= inputs(28);
    layer0_outputs(6818) <= (inputs(137)) or (inputs(87));
    layer0_outputs(6819) <= not((inputs(50)) or (inputs(86)));
    layer0_outputs(6820) <= not((inputs(198)) or (inputs(27)));
    layer0_outputs(6821) <= (inputs(112)) and not (inputs(206));
    layer0_outputs(6822) <= not((inputs(100)) xor (inputs(18)));
    layer0_outputs(6823) <= inputs(52);
    layer0_outputs(6824) <= not(inputs(73)) or (inputs(202));
    layer0_outputs(6825) <= (inputs(7)) xor (inputs(56));
    layer0_outputs(6826) <= (inputs(172)) and not (inputs(182));
    layer0_outputs(6827) <= not((inputs(22)) xor (inputs(85)));
    layer0_outputs(6828) <= (inputs(138)) and not (inputs(244));
    layer0_outputs(6829) <= not(inputs(167)) or (inputs(96));
    layer0_outputs(6830) <= not(inputs(21)) or (inputs(66));
    layer0_outputs(6831) <= not(inputs(82));
    layer0_outputs(6832) <= '0';
    layer0_outputs(6833) <= not(inputs(52));
    layer0_outputs(6834) <= not((inputs(91)) or (inputs(16)));
    layer0_outputs(6835) <= not(inputs(41));
    layer0_outputs(6836) <= not((inputs(21)) or (inputs(158)));
    layer0_outputs(6837) <= (inputs(36)) or (inputs(240));
    layer0_outputs(6838) <= (inputs(217)) or (inputs(28));
    layer0_outputs(6839) <= not((inputs(160)) xor (inputs(230)));
    layer0_outputs(6840) <= not((inputs(92)) and (inputs(92)));
    layer0_outputs(6841) <= (inputs(211)) and not (inputs(65));
    layer0_outputs(6842) <= not(inputs(159));
    layer0_outputs(6843) <= not(inputs(245));
    layer0_outputs(6844) <= inputs(97);
    layer0_outputs(6845) <= (inputs(18)) xor (inputs(180));
    layer0_outputs(6846) <= inputs(173);
    layer0_outputs(6847) <= '1';
    layer0_outputs(6848) <= not(inputs(114));
    layer0_outputs(6849) <= inputs(82);
    layer0_outputs(6850) <= inputs(120);
    layer0_outputs(6851) <= (inputs(125)) and not (inputs(225));
    layer0_outputs(6852) <= not(inputs(157)) or (inputs(32));
    layer0_outputs(6853) <= not(inputs(1));
    layer0_outputs(6854) <= not(inputs(141)) or (inputs(241));
    layer0_outputs(6855) <= not(inputs(189));
    layer0_outputs(6856) <= inputs(57);
    layer0_outputs(6857) <= (inputs(253)) or (inputs(143));
    layer0_outputs(6858) <= (inputs(55)) or (inputs(198));
    layer0_outputs(6859) <= not(inputs(221));
    layer0_outputs(6860) <= not(inputs(21)) or (inputs(208));
    layer0_outputs(6861) <= (inputs(208)) xor (inputs(184));
    layer0_outputs(6862) <= (inputs(120)) or (inputs(103));
    layer0_outputs(6863) <= not((inputs(218)) and (inputs(169)));
    layer0_outputs(6864) <= not((inputs(66)) or (inputs(195)));
    layer0_outputs(6865) <= not((inputs(218)) and (inputs(232)));
    layer0_outputs(6866) <= inputs(181);
    layer0_outputs(6867) <= (inputs(171)) or (inputs(100));
    layer0_outputs(6868) <= (inputs(189)) and not (inputs(162));
    layer0_outputs(6869) <= (inputs(110)) and (inputs(244));
    layer0_outputs(6870) <= (inputs(226)) or (inputs(134));
    layer0_outputs(6871) <= (inputs(233)) and not (inputs(3));
    layer0_outputs(6872) <= (inputs(233)) or (inputs(11));
    layer0_outputs(6873) <= not(inputs(177));
    layer0_outputs(6874) <= (inputs(79)) or (inputs(84));
    layer0_outputs(6875) <= not((inputs(39)) or (inputs(85)));
    layer0_outputs(6876) <= not(inputs(73)) or (inputs(251));
    layer0_outputs(6877) <= not(inputs(146));
    layer0_outputs(6878) <= not(inputs(49)) or (inputs(234));
    layer0_outputs(6879) <= not((inputs(239)) or (inputs(52)));
    layer0_outputs(6880) <= (inputs(25)) xor (inputs(113));
    layer0_outputs(6881) <= (inputs(68)) or (inputs(169));
    layer0_outputs(6882) <= (inputs(67)) or (inputs(85));
    layer0_outputs(6883) <= not((inputs(134)) or (inputs(165)));
    layer0_outputs(6884) <= not(inputs(215));
    layer0_outputs(6885) <= (inputs(66)) xor (inputs(77));
    layer0_outputs(6886) <= not((inputs(38)) xor (inputs(208)));
    layer0_outputs(6887) <= inputs(29);
    layer0_outputs(6888) <= (inputs(80)) xor (inputs(85));
    layer0_outputs(6889) <= not((inputs(14)) or (inputs(131)));
    layer0_outputs(6890) <= (inputs(190)) or (inputs(99));
    layer0_outputs(6891) <= not(inputs(23));
    layer0_outputs(6892) <= not(inputs(177)) or (inputs(224));
    layer0_outputs(6893) <= inputs(168);
    layer0_outputs(6894) <= not((inputs(123)) xor (inputs(155)));
    layer0_outputs(6895) <= inputs(9);
    layer0_outputs(6896) <= (inputs(8)) and not (inputs(239));
    layer0_outputs(6897) <= (inputs(245)) or (inputs(193));
    layer0_outputs(6898) <= (inputs(204)) or (inputs(220));
    layer0_outputs(6899) <= not((inputs(211)) and (inputs(11)));
    layer0_outputs(6900) <= not(inputs(114));
    layer0_outputs(6901) <= inputs(231);
    layer0_outputs(6902) <= (inputs(230)) and not (inputs(238));
    layer0_outputs(6903) <= not(inputs(223)) or (inputs(222));
    layer0_outputs(6904) <= inputs(108);
    layer0_outputs(6905) <= (inputs(58)) xor (inputs(11));
    layer0_outputs(6906) <= '1';
    layer0_outputs(6907) <= (inputs(216)) or (inputs(48));
    layer0_outputs(6908) <= not((inputs(5)) or (inputs(45)));
    layer0_outputs(6909) <= (inputs(207)) and not (inputs(187));
    layer0_outputs(6910) <= inputs(92);
    layer0_outputs(6911) <= (inputs(154)) and (inputs(55));
    layer0_outputs(6912) <= inputs(101);
    layer0_outputs(6913) <= (inputs(57)) or (inputs(13));
    layer0_outputs(6914) <= not(inputs(12));
    layer0_outputs(6915) <= not(inputs(237)) or (inputs(63));
    layer0_outputs(6916) <= not(inputs(239)) or (inputs(146));
    layer0_outputs(6917) <= not(inputs(173));
    layer0_outputs(6918) <= inputs(205);
    layer0_outputs(6919) <= inputs(180);
    layer0_outputs(6920) <= (inputs(138)) and not (inputs(233));
    layer0_outputs(6921) <= not(inputs(226));
    layer0_outputs(6922) <= (inputs(181)) or (inputs(108));
    layer0_outputs(6923) <= not(inputs(196));
    layer0_outputs(6924) <= '0';
    layer0_outputs(6925) <= not((inputs(75)) or (inputs(52)));
    layer0_outputs(6926) <= not((inputs(167)) xor (inputs(161)));
    layer0_outputs(6927) <= inputs(7);
    layer0_outputs(6928) <= not((inputs(87)) or (inputs(25)));
    layer0_outputs(6929) <= not(inputs(67)) or (inputs(50));
    layer0_outputs(6930) <= not(inputs(163)) or (inputs(176));
    layer0_outputs(6931) <= not(inputs(170)) or (inputs(153));
    layer0_outputs(6932) <= not((inputs(21)) xor (inputs(99)));
    layer0_outputs(6933) <= not((inputs(165)) and (inputs(217)));
    layer0_outputs(6934) <= (inputs(183)) or (inputs(87));
    layer0_outputs(6935) <= not(inputs(10));
    layer0_outputs(6936) <= inputs(215);
    layer0_outputs(6937) <= (inputs(59)) xor (inputs(61));
    layer0_outputs(6938) <= inputs(153);
    layer0_outputs(6939) <= '1';
    layer0_outputs(6940) <= not(inputs(230));
    layer0_outputs(6941) <= inputs(144);
    layer0_outputs(6942) <= inputs(142);
    layer0_outputs(6943) <= not((inputs(20)) or (inputs(174)));
    layer0_outputs(6944) <= not((inputs(138)) or (inputs(40)));
    layer0_outputs(6945) <= (inputs(125)) and not (inputs(254));
    layer0_outputs(6946) <= not(inputs(181));
    layer0_outputs(6947) <= not((inputs(166)) or (inputs(105)));
    layer0_outputs(6948) <= not(inputs(50));
    layer0_outputs(6949) <= not(inputs(89)) or (inputs(191));
    layer0_outputs(6950) <= not((inputs(172)) or (inputs(13)));
    layer0_outputs(6951) <= (inputs(246)) or (inputs(8));
    layer0_outputs(6952) <= (inputs(118)) xor (inputs(54));
    layer0_outputs(6953) <= not(inputs(132)) or (inputs(221));
    layer0_outputs(6954) <= not((inputs(208)) or (inputs(22)));
    layer0_outputs(6955) <= (inputs(59)) or (inputs(36));
    layer0_outputs(6956) <= inputs(169);
    layer0_outputs(6957) <= inputs(101);
    layer0_outputs(6958) <= '0';
    layer0_outputs(6959) <= inputs(24);
    layer0_outputs(6960) <= '1';
    layer0_outputs(6961) <= not((inputs(57)) and (inputs(7)));
    layer0_outputs(6962) <= not((inputs(157)) and (inputs(77)));
    layer0_outputs(6963) <= not((inputs(224)) xor (inputs(3)));
    layer0_outputs(6964) <= not((inputs(125)) or (inputs(126)));
    layer0_outputs(6965) <= not(inputs(248)) or (inputs(4));
    layer0_outputs(6966) <= (inputs(27)) and not (inputs(237));
    layer0_outputs(6967) <= not(inputs(57));
    layer0_outputs(6968) <= (inputs(142)) xor (inputs(122));
    layer0_outputs(6969) <= inputs(44);
    layer0_outputs(6970) <= (inputs(185)) and (inputs(187));
    layer0_outputs(6971) <= not(inputs(29)) or (inputs(186));
    layer0_outputs(6972) <= not((inputs(125)) and (inputs(229)));
    layer0_outputs(6973) <= (inputs(197)) or (inputs(141));
    layer0_outputs(6974) <= not(inputs(106));
    layer0_outputs(6975) <= not(inputs(160)) or (inputs(4));
    layer0_outputs(6976) <= (inputs(28)) and (inputs(28));
    layer0_outputs(6977) <= inputs(175);
    layer0_outputs(6978) <= not((inputs(18)) or (inputs(52)));
    layer0_outputs(6979) <= (inputs(75)) or (inputs(68));
    layer0_outputs(6980) <= (inputs(188)) or (inputs(173));
    layer0_outputs(6981) <= not(inputs(92));
    layer0_outputs(6982) <= (inputs(23)) and not (inputs(144));
    layer0_outputs(6983) <= (inputs(242)) xor (inputs(212));
    layer0_outputs(6984) <= not((inputs(186)) or (inputs(139)));
    layer0_outputs(6985) <= not((inputs(154)) or (inputs(222)));
    layer0_outputs(6986) <= not(inputs(125));
    layer0_outputs(6987) <= inputs(30);
    layer0_outputs(6988) <= not(inputs(239));
    layer0_outputs(6989) <= (inputs(241)) and not (inputs(244));
    layer0_outputs(6990) <= inputs(68);
    layer0_outputs(6991) <= (inputs(80)) and (inputs(194));
    layer0_outputs(6992) <= inputs(147);
    layer0_outputs(6993) <= (inputs(23)) or (inputs(207));
    layer0_outputs(6994) <= inputs(166);
    layer0_outputs(6995) <= not((inputs(17)) xor (inputs(132)));
    layer0_outputs(6996) <= not(inputs(162)) or (inputs(254));
    layer0_outputs(6997) <= (inputs(156)) or (inputs(243));
    layer0_outputs(6998) <= (inputs(254)) or (inputs(25));
    layer0_outputs(6999) <= not(inputs(133));
    layer0_outputs(7000) <= '0';
    layer0_outputs(7001) <= inputs(248);
    layer0_outputs(7002) <= inputs(230);
    layer0_outputs(7003) <= (inputs(194)) or (inputs(84));
    layer0_outputs(7004) <= (inputs(125)) and not (inputs(118));
    layer0_outputs(7005) <= (inputs(222)) xor (inputs(236));
    layer0_outputs(7006) <= inputs(203);
    layer0_outputs(7007) <= not(inputs(91)) or (inputs(214));
    layer0_outputs(7008) <= not(inputs(93)) or (inputs(184));
    layer0_outputs(7009) <= not((inputs(163)) and (inputs(55)));
    layer0_outputs(7010) <= inputs(52);
    layer0_outputs(7011) <= not(inputs(72)) or (inputs(80));
    layer0_outputs(7012) <= not(inputs(189)) or (inputs(55));
    layer0_outputs(7013) <= not(inputs(98));
    layer0_outputs(7014) <= inputs(89);
    layer0_outputs(7015) <= inputs(94);
    layer0_outputs(7016) <= (inputs(107)) xor (inputs(142));
    layer0_outputs(7017) <= inputs(71);
    layer0_outputs(7018) <= not(inputs(5));
    layer0_outputs(7019) <= '1';
    layer0_outputs(7020) <= not((inputs(212)) or (inputs(190)));
    layer0_outputs(7021) <= (inputs(76)) or (inputs(1));
    layer0_outputs(7022) <= not(inputs(138)) or (inputs(204));
    layer0_outputs(7023) <= (inputs(60)) or (inputs(137));
    layer0_outputs(7024) <= inputs(254);
    layer0_outputs(7025) <= (inputs(35)) or (inputs(91));
    layer0_outputs(7026) <= not((inputs(130)) xor (inputs(118)));
    layer0_outputs(7027) <= not(inputs(144)) or (inputs(174));
    layer0_outputs(7028) <= (inputs(8)) and (inputs(180));
    layer0_outputs(7029) <= (inputs(72)) or (inputs(126));
    layer0_outputs(7030) <= inputs(42);
    layer0_outputs(7031) <= not(inputs(114));
    layer0_outputs(7032) <= (inputs(74)) and not (inputs(41));
    layer0_outputs(7033) <= not((inputs(125)) or (inputs(176)));
    layer0_outputs(7034) <= not(inputs(145));
    layer0_outputs(7035) <= (inputs(253)) xor (inputs(161));
    layer0_outputs(7036) <= (inputs(23)) and not (inputs(250));
    layer0_outputs(7037) <= not(inputs(173));
    layer0_outputs(7038) <= (inputs(100)) xor (inputs(128));
    layer0_outputs(7039) <= inputs(196);
    layer0_outputs(7040) <= (inputs(190)) or (inputs(205));
    layer0_outputs(7041) <= (inputs(115)) or (inputs(82));
    layer0_outputs(7042) <= not((inputs(149)) and (inputs(230)));
    layer0_outputs(7043) <= (inputs(3)) xor (inputs(60));
    layer0_outputs(7044) <= not((inputs(234)) or (inputs(69)));
    layer0_outputs(7045) <= (inputs(237)) and not (inputs(190));
    layer0_outputs(7046) <= inputs(178);
    layer0_outputs(7047) <= not(inputs(84));
    layer0_outputs(7048) <= not(inputs(14));
    layer0_outputs(7049) <= (inputs(216)) or (inputs(113));
    layer0_outputs(7050) <= (inputs(177)) or (inputs(171));
    layer0_outputs(7051) <= '1';
    layer0_outputs(7052) <= not((inputs(38)) xor (inputs(159)));
    layer0_outputs(7053) <= inputs(123);
    layer0_outputs(7054) <= not((inputs(116)) xor (inputs(86)));
    layer0_outputs(7055) <= (inputs(52)) or (inputs(98));
    layer0_outputs(7056) <= (inputs(62)) or (inputs(246));
    layer0_outputs(7057) <= (inputs(242)) xor (inputs(58));
    layer0_outputs(7058) <= not(inputs(24));
    layer0_outputs(7059) <= inputs(163);
    layer0_outputs(7060) <= not(inputs(100));
    layer0_outputs(7061) <= not((inputs(21)) xor (inputs(57)));
    layer0_outputs(7062) <= inputs(62);
    layer0_outputs(7063) <= (inputs(125)) and not (inputs(128));
    layer0_outputs(7064) <= (inputs(6)) and not (inputs(130));
    layer0_outputs(7065) <= not(inputs(207));
    layer0_outputs(7066) <= (inputs(209)) or (inputs(49));
    layer0_outputs(7067) <= not((inputs(76)) xor (inputs(166)));
    layer0_outputs(7068) <= not(inputs(219));
    layer0_outputs(7069) <= (inputs(229)) or (inputs(205));
    layer0_outputs(7070) <= not(inputs(37));
    layer0_outputs(7071) <= (inputs(199)) xor (inputs(128));
    layer0_outputs(7072) <= (inputs(161)) or (inputs(76));
    layer0_outputs(7073) <= not(inputs(97)) or (inputs(157));
    layer0_outputs(7074) <= not(inputs(82)) or (inputs(106));
    layer0_outputs(7075) <= not(inputs(181));
    layer0_outputs(7076) <= not(inputs(135));
    layer0_outputs(7077) <= inputs(20);
    layer0_outputs(7078) <= inputs(98);
    layer0_outputs(7079) <= inputs(209);
    layer0_outputs(7080) <= not(inputs(198));
    layer0_outputs(7081) <= inputs(119);
    layer0_outputs(7082) <= (inputs(209)) or (inputs(41));
    layer0_outputs(7083) <= (inputs(63)) and not (inputs(95));
    layer0_outputs(7084) <= (inputs(172)) and not (inputs(99));
    layer0_outputs(7085) <= (inputs(90)) and not (inputs(177));
    layer0_outputs(7086) <= (inputs(0)) xor (inputs(90));
    layer0_outputs(7087) <= not(inputs(18));
    layer0_outputs(7088) <= (inputs(183)) or (inputs(177));
    layer0_outputs(7089) <= (inputs(128)) and not (inputs(135));
    layer0_outputs(7090) <= inputs(46);
    layer0_outputs(7091) <= (inputs(249)) or (inputs(180));
    layer0_outputs(7092) <= not((inputs(158)) xor (inputs(221)));
    layer0_outputs(7093) <= (inputs(196)) or (inputs(55));
    layer0_outputs(7094) <= not((inputs(7)) or (inputs(167)));
    layer0_outputs(7095) <= not((inputs(211)) or (inputs(87)));
    layer0_outputs(7096) <= inputs(24);
    layer0_outputs(7097) <= (inputs(184)) and (inputs(3));
    layer0_outputs(7098) <= not(inputs(228));
    layer0_outputs(7099) <= not(inputs(199)) or (inputs(141));
    layer0_outputs(7100) <= not(inputs(254)) or (inputs(58));
    layer0_outputs(7101) <= not(inputs(146));
    layer0_outputs(7102) <= '1';
    layer0_outputs(7103) <= not(inputs(197));
    layer0_outputs(7104) <= not(inputs(0)) or (inputs(205));
    layer0_outputs(7105) <= not(inputs(149));
    layer0_outputs(7106) <= not((inputs(171)) or (inputs(218)));
    layer0_outputs(7107) <= not((inputs(240)) and (inputs(0)));
    layer0_outputs(7108) <= not((inputs(25)) or (inputs(50)));
    layer0_outputs(7109) <= not((inputs(32)) and (inputs(120)));
    layer0_outputs(7110) <= (inputs(197)) or (inputs(116));
    layer0_outputs(7111) <= not((inputs(110)) or (inputs(153)));
    layer0_outputs(7112) <= inputs(198);
    layer0_outputs(7113) <= (inputs(221)) and not (inputs(157));
    layer0_outputs(7114) <= not(inputs(68)) or (inputs(126));
    layer0_outputs(7115) <= not((inputs(151)) or (inputs(237)));
    layer0_outputs(7116) <= '1';
    layer0_outputs(7117) <= not(inputs(113)) or (inputs(224));
    layer0_outputs(7118) <= not(inputs(75)) or (inputs(187));
    layer0_outputs(7119) <= (inputs(231)) and not (inputs(195));
    layer0_outputs(7120) <= inputs(23);
    layer0_outputs(7121) <= (inputs(227)) xor (inputs(207));
    layer0_outputs(7122) <= not((inputs(60)) or (inputs(230)));
    layer0_outputs(7123) <= (inputs(128)) and not (inputs(115));
    layer0_outputs(7124) <= inputs(188);
    layer0_outputs(7125) <= not((inputs(120)) and (inputs(89)));
    layer0_outputs(7126) <= (inputs(53)) xor (inputs(22));
    layer0_outputs(7127) <= not((inputs(254)) and (inputs(2)));
    layer0_outputs(7128) <= not(inputs(174));
    layer0_outputs(7129) <= not(inputs(220));
    layer0_outputs(7130) <= not(inputs(158));
    layer0_outputs(7131) <= not((inputs(80)) or (inputs(184)));
    layer0_outputs(7132) <= '0';
    layer0_outputs(7133) <= inputs(139);
    layer0_outputs(7134) <= not(inputs(87));
    layer0_outputs(7135) <= not(inputs(54));
    layer0_outputs(7136) <= not((inputs(54)) or (inputs(40)));
    layer0_outputs(7137) <= (inputs(68)) and not (inputs(62));
    layer0_outputs(7138) <= not((inputs(245)) and (inputs(217)));
    layer0_outputs(7139) <= (inputs(242)) or (inputs(11));
    layer0_outputs(7140) <= not((inputs(108)) or (inputs(164)));
    layer0_outputs(7141) <= not((inputs(146)) or (inputs(160)));
    layer0_outputs(7142) <= not(inputs(154)) or (inputs(212));
    layer0_outputs(7143) <= not(inputs(246));
    layer0_outputs(7144) <= inputs(169);
    layer0_outputs(7145) <= not(inputs(132));
    layer0_outputs(7146) <= (inputs(22)) or (inputs(67));
    layer0_outputs(7147) <= (inputs(145)) or (inputs(227));
    layer0_outputs(7148) <= (inputs(47)) or (inputs(153));
    layer0_outputs(7149) <= not(inputs(155)) or (inputs(16));
    layer0_outputs(7150) <= (inputs(161)) and not (inputs(53));
    layer0_outputs(7151) <= not(inputs(224)) or (inputs(16));
    layer0_outputs(7152) <= inputs(32);
    layer0_outputs(7153) <= not((inputs(142)) or (inputs(101)));
    layer0_outputs(7154) <= not(inputs(153));
    layer0_outputs(7155) <= (inputs(146)) and not (inputs(15));
    layer0_outputs(7156) <= (inputs(2)) or (inputs(202));
    layer0_outputs(7157) <= not(inputs(92));
    layer0_outputs(7158) <= (inputs(125)) and (inputs(185));
    layer0_outputs(7159) <= not((inputs(228)) or (inputs(67)));
    layer0_outputs(7160) <= '1';
    layer0_outputs(7161) <= (inputs(91)) or (inputs(12));
    layer0_outputs(7162) <= (inputs(16)) and not (inputs(114));
    layer0_outputs(7163) <= not((inputs(118)) or (inputs(100)));
    layer0_outputs(7164) <= not(inputs(65)) or (inputs(28));
    layer0_outputs(7165) <= not((inputs(119)) or (inputs(248)));
    layer0_outputs(7166) <= '0';
    layer0_outputs(7167) <= not(inputs(7)) or (inputs(84));
    layer0_outputs(7168) <= inputs(115);
    layer0_outputs(7169) <= (inputs(210)) and (inputs(70));
    layer0_outputs(7170) <= not((inputs(105)) or (inputs(93)));
    layer0_outputs(7171) <= not(inputs(107));
    layer0_outputs(7172) <= not((inputs(148)) xor (inputs(116)));
    layer0_outputs(7173) <= not(inputs(55)) or (inputs(56));
    layer0_outputs(7174) <= (inputs(226)) xor (inputs(206));
    layer0_outputs(7175) <= not((inputs(223)) or (inputs(161)));
    layer0_outputs(7176) <= inputs(196);
    layer0_outputs(7177) <= inputs(93);
    layer0_outputs(7178) <= (inputs(46)) or (inputs(169));
    layer0_outputs(7179) <= inputs(130);
    layer0_outputs(7180) <= (inputs(209)) or (inputs(125));
    layer0_outputs(7181) <= not(inputs(190));
    layer0_outputs(7182) <= not((inputs(215)) or (inputs(200)));
    layer0_outputs(7183) <= not(inputs(130));
    layer0_outputs(7184) <= (inputs(197)) and (inputs(159));
    layer0_outputs(7185) <= not(inputs(232));
    layer0_outputs(7186) <= not(inputs(187)) or (inputs(17));
    layer0_outputs(7187) <= inputs(101);
    layer0_outputs(7188) <= not((inputs(78)) or (inputs(210)));
    layer0_outputs(7189) <= not(inputs(24)) or (inputs(131));
    layer0_outputs(7190) <= (inputs(163)) and (inputs(255));
    layer0_outputs(7191) <= inputs(25);
    layer0_outputs(7192) <= not(inputs(145));
    layer0_outputs(7193) <= (inputs(210)) and (inputs(92));
    layer0_outputs(7194) <= inputs(23);
    layer0_outputs(7195) <= not((inputs(159)) and (inputs(111)));
    layer0_outputs(7196) <= inputs(180);
    layer0_outputs(7197) <= inputs(197);
    layer0_outputs(7198) <= not(inputs(167));
    layer0_outputs(7199) <= not(inputs(252));
    layer0_outputs(7200) <= (inputs(214)) or (inputs(205));
    layer0_outputs(7201) <= inputs(139);
    layer0_outputs(7202) <= (inputs(101)) and not (inputs(20));
    layer0_outputs(7203) <= not(inputs(91));
    layer0_outputs(7204) <= not((inputs(52)) xor (inputs(19)));
    layer0_outputs(7205) <= '1';
    layer0_outputs(7206) <= (inputs(1)) and not (inputs(41));
    layer0_outputs(7207) <= not((inputs(187)) or (inputs(242)));
    layer0_outputs(7208) <= inputs(66);
    layer0_outputs(7209) <= not(inputs(7)) or (inputs(163));
    layer0_outputs(7210) <= not((inputs(130)) or (inputs(5)));
    layer0_outputs(7211) <= inputs(226);
    layer0_outputs(7212) <= (inputs(36)) or (inputs(140));
    layer0_outputs(7213) <= not(inputs(124));
    layer0_outputs(7214) <= not(inputs(166)) or (inputs(184));
    layer0_outputs(7215) <= '1';
    layer0_outputs(7216) <= not((inputs(193)) or (inputs(19)));
    layer0_outputs(7217) <= (inputs(96)) or (inputs(146));
    layer0_outputs(7218) <= inputs(150);
    layer0_outputs(7219) <= not((inputs(86)) and (inputs(10)));
    layer0_outputs(7220) <= not((inputs(165)) xor (inputs(198)));
    layer0_outputs(7221) <= not(inputs(99)) or (inputs(200));
    layer0_outputs(7222) <= not((inputs(231)) and (inputs(228)));
    layer0_outputs(7223) <= inputs(168);
    layer0_outputs(7224) <= not((inputs(10)) xor (inputs(254)));
    layer0_outputs(7225) <= not(inputs(179));
    layer0_outputs(7226) <= inputs(179);
    layer0_outputs(7227) <= not(inputs(29)) or (inputs(45));
    layer0_outputs(7228) <= (inputs(2)) and not (inputs(254));
    layer0_outputs(7229) <= '1';
    layer0_outputs(7230) <= not((inputs(136)) and (inputs(196)));
    layer0_outputs(7231) <= not(inputs(102));
    layer0_outputs(7232) <= not((inputs(102)) xor (inputs(134)));
    layer0_outputs(7233) <= not(inputs(108));
    layer0_outputs(7234) <= not((inputs(83)) and (inputs(134)));
    layer0_outputs(7235) <= inputs(106);
    layer0_outputs(7236) <= (inputs(222)) and not (inputs(97));
    layer0_outputs(7237) <= not((inputs(154)) or (inputs(174)));
    layer0_outputs(7238) <= '0';
    layer0_outputs(7239) <= not((inputs(133)) or (inputs(179)));
    layer0_outputs(7240) <= (inputs(229)) and not (inputs(73));
    layer0_outputs(7241) <= not((inputs(99)) or (inputs(148)));
    layer0_outputs(7242) <= not((inputs(57)) or (inputs(159)));
    layer0_outputs(7243) <= not((inputs(136)) or (inputs(13)));
    layer0_outputs(7244) <= not(inputs(213)) or (inputs(59));
    layer0_outputs(7245) <= (inputs(110)) xor (inputs(208));
    layer0_outputs(7246) <= not(inputs(150)) or (inputs(84));
    layer0_outputs(7247) <= (inputs(240)) and not (inputs(51));
    layer0_outputs(7248) <= (inputs(43)) xor (inputs(175));
    layer0_outputs(7249) <= (inputs(81)) or (inputs(10));
    layer0_outputs(7250) <= '0';
    layer0_outputs(7251) <= (inputs(5)) xor (inputs(123));
    layer0_outputs(7252) <= (inputs(7)) and (inputs(211));
    layer0_outputs(7253) <= not((inputs(7)) or (inputs(4)));
    layer0_outputs(7254) <= not(inputs(98));
    layer0_outputs(7255) <= not((inputs(55)) or (inputs(75)));
    layer0_outputs(7256) <= inputs(33);
    layer0_outputs(7257) <= (inputs(16)) and (inputs(46));
    layer0_outputs(7258) <= not((inputs(227)) or (inputs(245)));
    layer0_outputs(7259) <= not(inputs(133)) or (inputs(251));
    layer0_outputs(7260) <= not(inputs(85));
    layer0_outputs(7261) <= not((inputs(110)) xor (inputs(194)));
    layer0_outputs(7262) <= not((inputs(34)) xor (inputs(252)));
    layer0_outputs(7263) <= not((inputs(74)) and (inputs(202)));
    layer0_outputs(7264) <= '0';
    layer0_outputs(7265) <= not(inputs(226));
    layer0_outputs(7266) <= not(inputs(121));
    layer0_outputs(7267) <= not((inputs(4)) and (inputs(0)));
    layer0_outputs(7268) <= not((inputs(246)) xor (inputs(192)));
    layer0_outputs(7269) <= not(inputs(235)) or (inputs(137));
    layer0_outputs(7270) <= not((inputs(57)) xor (inputs(181)));
    layer0_outputs(7271) <= not(inputs(217));
    layer0_outputs(7272) <= not(inputs(118)) or (inputs(4));
    layer0_outputs(7273) <= not((inputs(234)) or (inputs(48)));
    layer0_outputs(7274) <= (inputs(176)) and not (inputs(138));
    layer0_outputs(7275) <= not((inputs(108)) or (inputs(234)));
    layer0_outputs(7276) <= not((inputs(43)) or (inputs(110)));
    layer0_outputs(7277) <= (inputs(32)) and (inputs(169));
    layer0_outputs(7278) <= not((inputs(173)) xor (inputs(239)));
    layer0_outputs(7279) <= not((inputs(205)) or (inputs(182)));
    layer0_outputs(7280) <= inputs(252);
    layer0_outputs(7281) <= inputs(104);
    layer0_outputs(7282) <= (inputs(38)) and not (inputs(84));
    layer0_outputs(7283) <= (inputs(73)) and (inputs(130));
    layer0_outputs(7284) <= (inputs(138)) or (inputs(158));
    layer0_outputs(7285) <= inputs(121);
    layer0_outputs(7286) <= not((inputs(167)) or (inputs(201)));
    layer0_outputs(7287) <= not(inputs(103)) or (inputs(142));
    layer0_outputs(7288) <= not(inputs(28));
    layer0_outputs(7289) <= (inputs(171)) or (inputs(237));
    layer0_outputs(7290) <= (inputs(188)) and not (inputs(61));
    layer0_outputs(7291) <= (inputs(78)) and not (inputs(149));
    layer0_outputs(7292) <= (inputs(196)) and not (inputs(0));
    layer0_outputs(7293) <= not((inputs(65)) xor (inputs(103)));
    layer0_outputs(7294) <= not(inputs(237));
    layer0_outputs(7295) <= not((inputs(168)) or (inputs(20)));
    layer0_outputs(7296) <= (inputs(143)) or (inputs(126));
    layer0_outputs(7297) <= not((inputs(238)) or (inputs(220)));
    layer0_outputs(7298) <= (inputs(141)) and not (inputs(226));
    layer0_outputs(7299) <= inputs(114);
    layer0_outputs(7300) <= inputs(119);
    layer0_outputs(7301) <= (inputs(231)) and (inputs(114));
    layer0_outputs(7302) <= not(inputs(211)) or (inputs(182));
    layer0_outputs(7303) <= not(inputs(147)) or (inputs(33));
    layer0_outputs(7304) <= not(inputs(15));
    layer0_outputs(7305) <= '0';
    layer0_outputs(7306) <= '1';
    layer0_outputs(7307) <= not((inputs(48)) xor (inputs(172)));
    layer0_outputs(7308) <= inputs(87);
    layer0_outputs(7309) <= inputs(93);
    layer0_outputs(7310) <= not(inputs(156));
    layer0_outputs(7311) <= inputs(128);
    layer0_outputs(7312) <= not(inputs(135));
    layer0_outputs(7313) <= (inputs(22)) and not (inputs(186));
    layer0_outputs(7314) <= inputs(58);
    layer0_outputs(7315) <= '0';
    layer0_outputs(7316) <= (inputs(167)) or (inputs(226));
    layer0_outputs(7317) <= not((inputs(191)) and (inputs(82)));
    layer0_outputs(7318) <= '1';
    layer0_outputs(7319) <= not(inputs(195)) or (inputs(96));
    layer0_outputs(7320) <= (inputs(71)) and (inputs(28));
    layer0_outputs(7321) <= (inputs(148)) or (inputs(96));
    layer0_outputs(7322) <= inputs(155);
    layer0_outputs(7323) <= not(inputs(188));
    layer0_outputs(7324) <= not(inputs(208)) or (inputs(93));
    layer0_outputs(7325) <= not((inputs(17)) xor (inputs(199)));
    layer0_outputs(7326) <= not((inputs(170)) or (inputs(11)));
    layer0_outputs(7327) <= not((inputs(145)) or (inputs(232)));
    layer0_outputs(7328) <= not(inputs(157));
    layer0_outputs(7329) <= '0';
    layer0_outputs(7330) <= (inputs(147)) or (inputs(238));
    layer0_outputs(7331) <= not(inputs(102)) or (inputs(32));
    layer0_outputs(7332) <= not((inputs(128)) or (inputs(195)));
    layer0_outputs(7333) <= (inputs(120)) and not (inputs(253));
    layer0_outputs(7334) <= not(inputs(192));
    layer0_outputs(7335) <= not(inputs(135)) or (inputs(51));
    layer0_outputs(7336) <= (inputs(135)) and not (inputs(215));
    layer0_outputs(7337) <= (inputs(182)) or (inputs(5));
    layer0_outputs(7338) <= not((inputs(148)) or (inputs(180)));
    layer0_outputs(7339) <= (inputs(110)) and not (inputs(129));
    layer0_outputs(7340) <= (inputs(210)) and not (inputs(15));
    layer0_outputs(7341) <= inputs(114);
    layer0_outputs(7342) <= not(inputs(196)) or (inputs(133));
    layer0_outputs(7343) <= (inputs(154)) and not (inputs(14));
    layer0_outputs(7344) <= not(inputs(183));
    layer0_outputs(7345) <= not((inputs(85)) xor (inputs(23)));
    layer0_outputs(7346) <= inputs(135);
    layer0_outputs(7347) <= '0';
    layer0_outputs(7348) <= inputs(58);
    layer0_outputs(7349) <= not(inputs(7));
    layer0_outputs(7350) <= (inputs(23)) or (inputs(11));
    layer0_outputs(7351) <= (inputs(203)) xor (inputs(6));
    layer0_outputs(7352) <= inputs(229);
    layer0_outputs(7353) <= (inputs(238)) and not (inputs(61));
    layer0_outputs(7354) <= (inputs(247)) and not (inputs(214));
    layer0_outputs(7355) <= inputs(93);
    layer0_outputs(7356) <= (inputs(123)) and not (inputs(21));
    layer0_outputs(7357) <= not((inputs(30)) xor (inputs(29)));
    layer0_outputs(7358) <= (inputs(126)) or (inputs(78));
    layer0_outputs(7359) <= not(inputs(187));
    layer0_outputs(7360) <= not((inputs(236)) xor (inputs(191)));
    layer0_outputs(7361) <= '1';
    layer0_outputs(7362) <= (inputs(121)) and not (inputs(206));
    layer0_outputs(7363) <= not((inputs(78)) or (inputs(175)));
    layer0_outputs(7364) <= '1';
    layer0_outputs(7365) <= not(inputs(75));
    layer0_outputs(7366) <= (inputs(132)) and not (inputs(55));
    layer0_outputs(7367) <= '0';
    layer0_outputs(7368) <= (inputs(135)) or (inputs(166));
    layer0_outputs(7369) <= (inputs(132)) or (inputs(17));
    layer0_outputs(7370) <= inputs(24);
    layer0_outputs(7371) <= not(inputs(85));
    layer0_outputs(7372) <= inputs(5);
    layer0_outputs(7373) <= not(inputs(220));
    layer0_outputs(7374) <= not((inputs(128)) or (inputs(35)));
    layer0_outputs(7375) <= (inputs(242)) and not (inputs(242));
    layer0_outputs(7376) <= (inputs(105)) and not (inputs(126));
    layer0_outputs(7377) <= not(inputs(148));
    layer0_outputs(7378) <= (inputs(124)) and not (inputs(211));
    layer0_outputs(7379) <= not((inputs(247)) and (inputs(36)));
    layer0_outputs(7380) <= not((inputs(50)) xor (inputs(132)));
    layer0_outputs(7381) <= not(inputs(233));
    layer0_outputs(7382) <= (inputs(63)) and not (inputs(50));
    layer0_outputs(7383) <= not(inputs(19)) or (inputs(248));
    layer0_outputs(7384) <= not(inputs(232));
    layer0_outputs(7385) <= inputs(123);
    layer0_outputs(7386) <= not((inputs(135)) and (inputs(90)));
    layer0_outputs(7387) <= (inputs(95)) and not (inputs(123));
    layer0_outputs(7388) <= not(inputs(231));
    layer0_outputs(7389) <= (inputs(247)) or (inputs(187));
    layer0_outputs(7390) <= inputs(107);
    layer0_outputs(7391) <= not(inputs(190)) or (inputs(7));
    layer0_outputs(7392) <= (inputs(112)) or (inputs(65));
    layer0_outputs(7393) <= not(inputs(109));
    layer0_outputs(7394) <= not((inputs(32)) or (inputs(141)));
    layer0_outputs(7395) <= (inputs(222)) or (inputs(184));
    layer0_outputs(7396) <= inputs(10);
    layer0_outputs(7397) <= not(inputs(193));
    layer0_outputs(7398) <= not(inputs(84));
    layer0_outputs(7399) <= not((inputs(152)) and (inputs(217)));
    layer0_outputs(7400) <= inputs(181);
    layer0_outputs(7401) <= not((inputs(155)) xor (inputs(229)));
    layer0_outputs(7402) <= (inputs(61)) and not (inputs(128));
    layer0_outputs(7403) <= not((inputs(19)) or (inputs(31)));
    layer0_outputs(7404) <= inputs(90);
    layer0_outputs(7405) <= not(inputs(76));
    layer0_outputs(7406) <= (inputs(5)) or (inputs(143));
    layer0_outputs(7407) <= not((inputs(177)) or (inputs(246)));
    layer0_outputs(7408) <= not((inputs(236)) or (inputs(183)));
    layer0_outputs(7409) <= (inputs(73)) and not (inputs(182));
    layer0_outputs(7410) <= inputs(214);
    layer0_outputs(7411) <= not((inputs(187)) and (inputs(40)));
    layer0_outputs(7412) <= (inputs(31)) xor (inputs(116));
    layer0_outputs(7413) <= not(inputs(137));
    layer0_outputs(7414) <= not(inputs(234));
    layer0_outputs(7415) <= '0';
    layer0_outputs(7416) <= not(inputs(36));
    layer0_outputs(7417) <= (inputs(100)) or (inputs(83));
    layer0_outputs(7418) <= (inputs(81)) xor (inputs(67));
    layer0_outputs(7419) <= (inputs(189)) or (inputs(124));
    layer0_outputs(7420) <= not((inputs(113)) and (inputs(96)));
    layer0_outputs(7421) <= not(inputs(59));
    layer0_outputs(7422) <= inputs(210);
    layer0_outputs(7423) <= not((inputs(19)) or (inputs(215)));
    layer0_outputs(7424) <= (inputs(211)) or (inputs(243));
    layer0_outputs(7425) <= not(inputs(101)) or (inputs(181));
    layer0_outputs(7426) <= inputs(162);
    layer0_outputs(7427) <= inputs(141);
    layer0_outputs(7428) <= not(inputs(150));
    layer0_outputs(7429) <= not(inputs(244)) or (inputs(96));
    layer0_outputs(7430) <= '1';
    layer0_outputs(7431) <= not((inputs(75)) or (inputs(33)));
    layer0_outputs(7432) <= (inputs(153)) xor (inputs(30));
    layer0_outputs(7433) <= not((inputs(108)) or (inputs(187)));
    layer0_outputs(7434) <= not(inputs(228)) or (inputs(2));
    layer0_outputs(7435) <= not(inputs(48)) or (inputs(249));
    layer0_outputs(7436) <= (inputs(47)) and not (inputs(164));
    layer0_outputs(7437) <= not((inputs(235)) and (inputs(193)));
    layer0_outputs(7438) <= not((inputs(130)) or (inputs(100)));
    layer0_outputs(7439) <= not(inputs(218)) or (inputs(97));
    layer0_outputs(7440) <= not((inputs(228)) and (inputs(181)));
    layer0_outputs(7441) <= not((inputs(47)) or (inputs(73)));
    layer0_outputs(7442) <= '0';
    layer0_outputs(7443) <= (inputs(222)) or (inputs(76));
    layer0_outputs(7444) <= inputs(66);
    layer0_outputs(7445) <= (inputs(67)) or (inputs(80));
    layer0_outputs(7446) <= not(inputs(41));
    layer0_outputs(7447) <= inputs(255);
    layer0_outputs(7448) <= inputs(137);
    layer0_outputs(7449) <= (inputs(203)) or (inputs(156));
    layer0_outputs(7450) <= inputs(166);
    layer0_outputs(7451) <= (inputs(57)) and not (inputs(83));
    layer0_outputs(7452) <= inputs(39);
    layer0_outputs(7453) <= not(inputs(208));
    layer0_outputs(7454) <= (inputs(192)) or (inputs(126));
    layer0_outputs(7455) <= (inputs(131)) or (inputs(247));
    layer0_outputs(7456) <= (inputs(19)) or (inputs(32));
    layer0_outputs(7457) <= (inputs(75)) and not (inputs(47));
    layer0_outputs(7458) <= (inputs(96)) or (inputs(191));
    layer0_outputs(7459) <= (inputs(86)) or (inputs(203));
    layer0_outputs(7460) <= (inputs(118)) or (inputs(104));
    layer0_outputs(7461) <= not(inputs(223)) or (inputs(49));
    layer0_outputs(7462) <= (inputs(218)) and not (inputs(231));
    layer0_outputs(7463) <= (inputs(197)) xor (inputs(59));
    layer0_outputs(7464) <= not((inputs(6)) or (inputs(13)));
    layer0_outputs(7465) <= inputs(39);
    layer0_outputs(7466) <= inputs(115);
    layer0_outputs(7467) <= not((inputs(191)) or (inputs(55)));
    layer0_outputs(7468) <= not((inputs(168)) xor (inputs(64)));
    layer0_outputs(7469) <= inputs(204);
    layer0_outputs(7470) <= not(inputs(114));
    layer0_outputs(7471) <= not(inputs(112));
    layer0_outputs(7472) <= '0';
    layer0_outputs(7473) <= not((inputs(46)) or (inputs(38)));
    layer0_outputs(7474) <= inputs(21);
    layer0_outputs(7475) <= inputs(149);
    layer0_outputs(7476) <= (inputs(242)) and not (inputs(31));
    layer0_outputs(7477) <= not(inputs(130));
    layer0_outputs(7478) <= inputs(161);
    layer0_outputs(7479) <= not((inputs(82)) or (inputs(79)));
    layer0_outputs(7480) <= not(inputs(120));
    layer0_outputs(7481) <= not(inputs(182));
    layer0_outputs(7482) <= not(inputs(68)) or (inputs(73));
    layer0_outputs(7483) <= inputs(62);
    layer0_outputs(7484) <= not((inputs(67)) xor (inputs(53)));
    layer0_outputs(7485) <= inputs(199);
    layer0_outputs(7486) <= not((inputs(75)) xor (inputs(59)));
    layer0_outputs(7487) <= inputs(94);
    layer0_outputs(7488) <= not((inputs(130)) xor (inputs(181)));
    layer0_outputs(7489) <= not(inputs(113)) or (inputs(139));
    layer0_outputs(7490) <= inputs(109);
    layer0_outputs(7491) <= not(inputs(100)) or (inputs(8));
    layer0_outputs(7492) <= (inputs(105)) or (inputs(79));
    layer0_outputs(7493) <= not((inputs(130)) xor (inputs(183)));
    layer0_outputs(7494) <= not((inputs(196)) or (inputs(146)));
    layer0_outputs(7495) <= not((inputs(55)) or (inputs(220)));
    layer0_outputs(7496) <= not(inputs(103)) or (inputs(162));
    layer0_outputs(7497) <= (inputs(202)) or (inputs(88));
    layer0_outputs(7498) <= not(inputs(245)) or (inputs(36));
    layer0_outputs(7499) <= not((inputs(157)) or (inputs(156)));
    layer0_outputs(7500) <= not((inputs(217)) or (inputs(190)));
    layer0_outputs(7501) <= not(inputs(109)) or (inputs(89));
    layer0_outputs(7502) <= not(inputs(121));
    layer0_outputs(7503) <= (inputs(110)) or (inputs(251));
    layer0_outputs(7504) <= not(inputs(62));
    layer0_outputs(7505) <= (inputs(204)) or (inputs(58));
    layer0_outputs(7506) <= inputs(131);
    layer0_outputs(7507) <= (inputs(85)) xor (inputs(53));
    layer0_outputs(7508) <= not(inputs(233));
    layer0_outputs(7509) <= inputs(169);
    layer0_outputs(7510) <= not((inputs(197)) or (inputs(220)));
    layer0_outputs(7511) <= not(inputs(37));
    layer0_outputs(7512) <= inputs(121);
    layer0_outputs(7513) <= (inputs(245)) and not (inputs(236));
    layer0_outputs(7514) <= (inputs(23)) and not (inputs(96));
    layer0_outputs(7515) <= '1';
    layer0_outputs(7516) <= inputs(90);
    layer0_outputs(7517) <= (inputs(235)) and not (inputs(125));
    layer0_outputs(7518) <= not((inputs(71)) and (inputs(56)));
    layer0_outputs(7519) <= not(inputs(186));
    layer0_outputs(7520) <= '0';
    layer0_outputs(7521) <= inputs(156);
    layer0_outputs(7522) <= (inputs(149)) and not (inputs(13));
    layer0_outputs(7523) <= '1';
    layer0_outputs(7524) <= not(inputs(61));
    layer0_outputs(7525) <= inputs(250);
    layer0_outputs(7526) <= not(inputs(105)) or (inputs(180));
    layer0_outputs(7527) <= not(inputs(165)) or (inputs(132));
    layer0_outputs(7528) <= (inputs(44)) and not (inputs(105));
    layer0_outputs(7529) <= (inputs(108)) or (inputs(30));
    layer0_outputs(7530) <= (inputs(112)) and not (inputs(85));
    layer0_outputs(7531) <= inputs(145);
    layer0_outputs(7532) <= (inputs(68)) and (inputs(247));
    layer0_outputs(7533) <= not(inputs(36)) or (inputs(221));
    layer0_outputs(7534) <= not((inputs(212)) and (inputs(201)));
    layer0_outputs(7535) <= (inputs(8)) and not (inputs(2));
    layer0_outputs(7536) <= not(inputs(220));
    layer0_outputs(7537) <= '1';
    layer0_outputs(7538) <= not((inputs(37)) or (inputs(248)));
    layer0_outputs(7539) <= not(inputs(251));
    layer0_outputs(7540) <= '1';
    layer0_outputs(7541) <= not(inputs(94));
    layer0_outputs(7542) <= inputs(2);
    layer0_outputs(7543) <= (inputs(163)) or (inputs(142));
    layer0_outputs(7544) <= '0';
    layer0_outputs(7545) <= inputs(153);
    layer0_outputs(7546) <= not(inputs(132));
    layer0_outputs(7547) <= (inputs(205)) or (inputs(149));
    layer0_outputs(7548) <= not(inputs(219)) or (inputs(200));
    layer0_outputs(7549) <= (inputs(146)) or (inputs(202));
    layer0_outputs(7550) <= not(inputs(189)) or (inputs(162));
    layer0_outputs(7551) <= (inputs(153)) xor (inputs(32));
    layer0_outputs(7552) <= (inputs(145)) and not (inputs(255));
    layer0_outputs(7553) <= not((inputs(153)) and (inputs(202)));
    layer0_outputs(7554) <= (inputs(162)) and not (inputs(15));
    layer0_outputs(7555) <= (inputs(122)) and not (inputs(228));
    layer0_outputs(7556) <= inputs(179);
    layer0_outputs(7557) <= (inputs(6)) xor (inputs(199));
    layer0_outputs(7558) <= not((inputs(229)) and (inputs(104)));
    layer0_outputs(7559) <= (inputs(36)) and not (inputs(237));
    layer0_outputs(7560) <= not(inputs(65));
    layer0_outputs(7561) <= not((inputs(149)) or (inputs(122)));
    layer0_outputs(7562) <= not(inputs(119));
    layer0_outputs(7563) <= (inputs(88)) or (inputs(220));
    layer0_outputs(7564) <= not(inputs(164)) or (inputs(51));
    layer0_outputs(7565) <= not((inputs(194)) and (inputs(70)));
    layer0_outputs(7566) <= not(inputs(138)) or (inputs(237));
    layer0_outputs(7567) <= (inputs(241)) and not (inputs(159));
    layer0_outputs(7568) <= inputs(183);
    layer0_outputs(7569) <= (inputs(21)) and not (inputs(225));
    layer0_outputs(7570) <= inputs(111);
    layer0_outputs(7571) <= not(inputs(201)) or (inputs(83));
    layer0_outputs(7572) <= not(inputs(228));
    layer0_outputs(7573) <= not(inputs(0));
    layer0_outputs(7574) <= (inputs(28)) and not (inputs(171));
    layer0_outputs(7575) <= (inputs(171)) and not (inputs(52));
    layer0_outputs(7576) <= not(inputs(245));
    layer0_outputs(7577) <= not(inputs(165));
    layer0_outputs(7578) <= (inputs(183)) and (inputs(241));
    layer0_outputs(7579) <= (inputs(186)) and not (inputs(121));
    layer0_outputs(7580) <= not(inputs(9)) or (inputs(159));
    layer0_outputs(7581) <= (inputs(21)) or (inputs(124));
    layer0_outputs(7582) <= inputs(196);
    layer0_outputs(7583) <= (inputs(1)) or (inputs(59));
    layer0_outputs(7584) <= (inputs(37)) and not (inputs(144));
    layer0_outputs(7585) <= '0';
    layer0_outputs(7586) <= (inputs(252)) xor (inputs(203));
    layer0_outputs(7587) <= not(inputs(49));
    layer0_outputs(7588) <= (inputs(145)) xor (inputs(73));
    layer0_outputs(7589) <= not((inputs(80)) or (inputs(247)));
    layer0_outputs(7590) <= not((inputs(245)) or (inputs(62)));
    layer0_outputs(7591) <= inputs(159);
    layer0_outputs(7592) <= not(inputs(227)) or (inputs(112));
    layer0_outputs(7593) <= not(inputs(67));
    layer0_outputs(7594) <= inputs(119);
    layer0_outputs(7595) <= not((inputs(21)) and (inputs(92)));
    layer0_outputs(7596) <= not((inputs(96)) or (inputs(79)));
    layer0_outputs(7597) <= (inputs(167)) and not (inputs(105));
    layer0_outputs(7598) <= not((inputs(75)) or (inputs(11)));
    layer0_outputs(7599) <= not(inputs(42)) or (inputs(102));
    layer0_outputs(7600) <= inputs(119);
    layer0_outputs(7601) <= not((inputs(238)) or (inputs(159)));
    layer0_outputs(7602) <= inputs(229);
    layer0_outputs(7603) <= not((inputs(104)) or (inputs(138)));
    layer0_outputs(7604) <= not(inputs(77));
    layer0_outputs(7605) <= (inputs(31)) and (inputs(15));
    layer0_outputs(7606) <= not(inputs(17)) or (inputs(245));
    layer0_outputs(7607) <= not(inputs(87));
    layer0_outputs(7608) <= not((inputs(176)) or (inputs(208)));
    layer0_outputs(7609) <= (inputs(72)) or (inputs(250));
    layer0_outputs(7610) <= (inputs(105)) and not (inputs(228));
    layer0_outputs(7611) <= not(inputs(92));
    layer0_outputs(7612) <= (inputs(208)) and not (inputs(47));
    layer0_outputs(7613) <= not((inputs(61)) or (inputs(106)));
    layer0_outputs(7614) <= not((inputs(156)) or (inputs(234)));
    layer0_outputs(7615) <= not(inputs(179)) or (inputs(13));
    layer0_outputs(7616) <= not(inputs(38)) or (inputs(99));
    layer0_outputs(7617) <= '0';
    layer0_outputs(7618) <= inputs(104);
    layer0_outputs(7619) <= inputs(84);
    layer0_outputs(7620) <= (inputs(4)) and not (inputs(112));
    layer0_outputs(7621) <= inputs(15);
    layer0_outputs(7622) <= not((inputs(217)) or (inputs(207)));
    layer0_outputs(7623) <= (inputs(138)) and not (inputs(144));
    layer0_outputs(7624) <= inputs(214);
    layer0_outputs(7625) <= '1';
    layer0_outputs(7626) <= (inputs(54)) or (inputs(3));
    layer0_outputs(7627) <= not(inputs(92));
    layer0_outputs(7628) <= inputs(38);
    layer0_outputs(7629) <= (inputs(186)) or (inputs(4));
    layer0_outputs(7630) <= '1';
    layer0_outputs(7631) <= not(inputs(122));
    layer0_outputs(7632) <= not(inputs(82));
    layer0_outputs(7633) <= not((inputs(41)) and (inputs(214)));
    layer0_outputs(7634) <= inputs(132);
    layer0_outputs(7635) <= not(inputs(25)) or (inputs(40));
    layer0_outputs(7636) <= (inputs(239)) xor (inputs(104));
    layer0_outputs(7637) <= not((inputs(109)) or (inputs(85)));
    layer0_outputs(7638) <= inputs(204);
    layer0_outputs(7639) <= not((inputs(244)) or (inputs(5)));
    layer0_outputs(7640) <= (inputs(231)) and not (inputs(148));
    layer0_outputs(7641) <= '0';
    layer0_outputs(7642) <= (inputs(179)) and not (inputs(97));
    layer0_outputs(7643) <= not(inputs(178));
    layer0_outputs(7644) <= inputs(135);
    layer0_outputs(7645) <= inputs(26);
    layer0_outputs(7646) <= (inputs(112)) and (inputs(7));
    layer0_outputs(7647) <= inputs(254);
    layer0_outputs(7648) <= inputs(101);
    layer0_outputs(7649) <= (inputs(63)) and not (inputs(156));
    layer0_outputs(7650) <= '0';
    layer0_outputs(7651) <= not(inputs(26));
    layer0_outputs(7652) <= inputs(98);
    layer0_outputs(7653) <= (inputs(4)) and (inputs(90));
    layer0_outputs(7654) <= not((inputs(15)) or (inputs(108)));
    layer0_outputs(7655) <= not(inputs(183));
    layer0_outputs(7656) <= not((inputs(26)) or (inputs(233)));
    layer0_outputs(7657) <= not(inputs(90)) or (inputs(145));
    layer0_outputs(7658) <= not(inputs(162));
    layer0_outputs(7659) <= (inputs(153)) and (inputs(249));
    layer0_outputs(7660) <= not(inputs(221));
    layer0_outputs(7661) <= (inputs(19)) xor (inputs(39));
    layer0_outputs(7662) <= (inputs(73)) and not (inputs(49));
    layer0_outputs(7663) <= (inputs(51)) xor (inputs(46));
    layer0_outputs(7664) <= inputs(169);
    layer0_outputs(7665) <= (inputs(136)) xor (inputs(111));
    layer0_outputs(7666) <= (inputs(174)) xor (inputs(170));
    layer0_outputs(7667) <= not(inputs(71));
    layer0_outputs(7668) <= not((inputs(140)) xor (inputs(82)));
    layer0_outputs(7669) <= '1';
    layer0_outputs(7670) <= not((inputs(104)) or (inputs(20)));
    layer0_outputs(7671) <= not(inputs(84));
    layer0_outputs(7672) <= not((inputs(85)) or (inputs(127)));
    layer0_outputs(7673) <= not((inputs(18)) or (inputs(34)));
    layer0_outputs(7674) <= not(inputs(193)) or (inputs(157));
    layer0_outputs(7675) <= (inputs(72)) and (inputs(21));
    layer0_outputs(7676) <= (inputs(226)) and not (inputs(61));
    layer0_outputs(7677) <= not((inputs(142)) xor (inputs(197)));
    layer0_outputs(7678) <= not((inputs(234)) or (inputs(88)));
    layer0_outputs(7679) <= inputs(118);
    layer0_outputs(7680) <= not((inputs(22)) xor (inputs(27)));
    layer0_outputs(7681) <= not((inputs(50)) or (inputs(151)));
    layer0_outputs(7682) <= not((inputs(171)) or (inputs(248)));
    layer0_outputs(7683) <= (inputs(13)) or (inputs(120));
    layer0_outputs(7684) <= (inputs(164)) and not (inputs(83));
    layer0_outputs(7685) <= not((inputs(112)) or (inputs(17)));
    layer0_outputs(7686) <= (inputs(79)) xor (inputs(188));
    layer0_outputs(7687) <= '1';
    layer0_outputs(7688) <= (inputs(111)) or (inputs(51));
    layer0_outputs(7689) <= not(inputs(122)) or (inputs(47));
    layer0_outputs(7690) <= not((inputs(240)) and (inputs(194)));
    layer0_outputs(7691) <= not((inputs(126)) and (inputs(58)));
    layer0_outputs(7692) <= inputs(100);
    layer0_outputs(7693) <= inputs(117);
    layer0_outputs(7694) <= (inputs(34)) and (inputs(42));
    layer0_outputs(7695) <= not((inputs(0)) and (inputs(169)));
    layer0_outputs(7696) <= inputs(11);
    layer0_outputs(7697) <= (inputs(42)) and not (inputs(3));
    layer0_outputs(7698) <= not(inputs(55)) or (inputs(80));
    layer0_outputs(7699) <= (inputs(255)) and not (inputs(170));
    layer0_outputs(7700) <= (inputs(142)) and (inputs(198));
    layer0_outputs(7701) <= inputs(209);
    layer0_outputs(7702) <= inputs(102);
    layer0_outputs(7703) <= (inputs(58)) and not (inputs(165));
    layer0_outputs(7704) <= inputs(25);
    layer0_outputs(7705) <= inputs(167);
    layer0_outputs(7706) <= not((inputs(243)) or (inputs(153)));
    layer0_outputs(7707) <= inputs(72);
    layer0_outputs(7708) <= (inputs(231)) and not (inputs(7));
    layer0_outputs(7709) <= inputs(40);
    layer0_outputs(7710) <= (inputs(20)) and not (inputs(135));
    layer0_outputs(7711) <= inputs(25);
    layer0_outputs(7712) <= (inputs(181)) or (inputs(237));
    layer0_outputs(7713) <= inputs(136);
    layer0_outputs(7714) <= (inputs(54)) xor (inputs(79));
    layer0_outputs(7715) <= (inputs(67)) xor (inputs(190));
    layer0_outputs(7716) <= inputs(220);
    layer0_outputs(7717) <= inputs(60);
    layer0_outputs(7718) <= not((inputs(195)) and (inputs(212)));
    layer0_outputs(7719) <= inputs(27);
    layer0_outputs(7720) <= not((inputs(191)) or (inputs(144)));
    layer0_outputs(7721) <= not((inputs(178)) or (inputs(223)));
    layer0_outputs(7722) <= not((inputs(124)) and (inputs(44)));
    layer0_outputs(7723) <= not(inputs(131));
    layer0_outputs(7724) <= not(inputs(100));
    layer0_outputs(7725) <= inputs(254);
    layer0_outputs(7726) <= (inputs(233)) and (inputs(138));
    layer0_outputs(7727) <= (inputs(220)) xor (inputs(172));
    layer0_outputs(7728) <= not((inputs(48)) or (inputs(41)));
    layer0_outputs(7729) <= (inputs(79)) or (inputs(25));
    layer0_outputs(7730) <= inputs(119);
    layer0_outputs(7731) <= '0';
    layer0_outputs(7732) <= (inputs(66)) xor (inputs(231));
    layer0_outputs(7733) <= not((inputs(22)) or (inputs(31)));
    layer0_outputs(7734) <= not(inputs(132));
    layer0_outputs(7735) <= not(inputs(111));
    layer0_outputs(7736) <= not(inputs(142));
    layer0_outputs(7737) <= not(inputs(84));
    layer0_outputs(7738) <= (inputs(175)) and not (inputs(58));
    layer0_outputs(7739) <= (inputs(46)) and (inputs(108));
    layer0_outputs(7740) <= '0';
    layer0_outputs(7741) <= (inputs(226)) or (inputs(237));
    layer0_outputs(7742) <= not((inputs(142)) xor (inputs(94)));
    layer0_outputs(7743) <= inputs(46);
    layer0_outputs(7744) <= inputs(149);
    layer0_outputs(7745) <= not(inputs(128)) or (inputs(80));
    layer0_outputs(7746) <= inputs(20);
    layer0_outputs(7747) <= not(inputs(100)) or (inputs(251));
    layer0_outputs(7748) <= not(inputs(41)) or (inputs(1));
    layer0_outputs(7749) <= not(inputs(154)) or (inputs(186));
    layer0_outputs(7750) <= '0';
    layer0_outputs(7751) <= not((inputs(60)) or (inputs(46)));
    layer0_outputs(7752) <= (inputs(39)) and not (inputs(15));
    layer0_outputs(7753) <= not((inputs(171)) or (inputs(163)));
    layer0_outputs(7754) <= not((inputs(13)) or (inputs(16)));
    layer0_outputs(7755) <= '0';
    layer0_outputs(7756) <= not((inputs(108)) or (inputs(147)));
    layer0_outputs(7757) <= '0';
    layer0_outputs(7758) <= (inputs(158)) or (inputs(193));
    layer0_outputs(7759) <= (inputs(3)) and (inputs(39));
    layer0_outputs(7760) <= not((inputs(160)) or (inputs(144)));
    layer0_outputs(7761) <= not((inputs(233)) and (inputs(173)));
    layer0_outputs(7762) <= not(inputs(155));
    layer0_outputs(7763) <= '0';
    layer0_outputs(7764) <= not((inputs(202)) or (inputs(208)));
    layer0_outputs(7765) <= not(inputs(190));
    layer0_outputs(7766) <= (inputs(78)) xor (inputs(19));
    layer0_outputs(7767) <= not(inputs(22)) or (inputs(111));
    layer0_outputs(7768) <= not((inputs(125)) or (inputs(43)));
    layer0_outputs(7769) <= inputs(108);
    layer0_outputs(7770) <= inputs(225);
    layer0_outputs(7771) <= '1';
    layer0_outputs(7772) <= not((inputs(239)) xor (inputs(248)));
    layer0_outputs(7773) <= (inputs(71)) xor (inputs(16));
    layer0_outputs(7774) <= not((inputs(101)) or (inputs(29)));
    layer0_outputs(7775) <= not((inputs(250)) or (inputs(248)));
    layer0_outputs(7776) <= inputs(83);
    layer0_outputs(7777) <= inputs(219);
    layer0_outputs(7778) <= inputs(163);
    layer0_outputs(7779) <= (inputs(207)) and (inputs(108));
    layer0_outputs(7780) <= (inputs(29)) and (inputs(142));
    layer0_outputs(7781) <= (inputs(107)) or (inputs(4));
    layer0_outputs(7782) <= '1';
    layer0_outputs(7783) <= '0';
    layer0_outputs(7784) <= inputs(162);
    layer0_outputs(7785) <= not(inputs(28)) or (inputs(205));
    layer0_outputs(7786) <= not(inputs(26));
    layer0_outputs(7787) <= '0';
    layer0_outputs(7788) <= (inputs(217)) and not (inputs(121));
    layer0_outputs(7789) <= not(inputs(89)) or (inputs(124));
    layer0_outputs(7790) <= inputs(216);
    layer0_outputs(7791) <= not((inputs(194)) or (inputs(191)));
    layer0_outputs(7792) <= not((inputs(164)) xor (inputs(146)));
    layer0_outputs(7793) <= not((inputs(27)) or (inputs(214)));
    layer0_outputs(7794) <= inputs(151);
    layer0_outputs(7795) <= inputs(73);
    layer0_outputs(7796) <= (inputs(202)) or (inputs(141));
    layer0_outputs(7797) <= not(inputs(173));
    layer0_outputs(7798) <= not(inputs(133));
    layer0_outputs(7799) <= (inputs(159)) and not (inputs(137));
    layer0_outputs(7800) <= not(inputs(224)) or (inputs(0));
    layer0_outputs(7801) <= inputs(148);
    layer0_outputs(7802) <= (inputs(149)) and not (inputs(136));
    layer0_outputs(7803) <= not(inputs(140)) or (inputs(198));
    layer0_outputs(7804) <= not(inputs(40)) or (inputs(31));
    layer0_outputs(7805) <= not((inputs(6)) or (inputs(91)));
    layer0_outputs(7806) <= inputs(153);
    layer0_outputs(7807) <= (inputs(172)) and not (inputs(81));
    layer0_outputs(7808) <= inputs(38);
    layer0_outputs(7809) <= not((inputs(249)) xor (inputs(177)));
    layer0_outputs(7810) <= (inputs(37)) and not (inputs(129));
    layer0_outputs(7811) <= (inputs(148)) and (inputs(72));
    layer0_outputs(7812) <= inputs(221);
    layer0_outputs(7813) <= '0';
    layer0_outputs(7814) <= (inputs(10)) and not (inputs(184));
    layer0_outputs(7815) <= not(inputs(139));
    layer0_outputs(7816) <= (inputs(98)) or (inputs(247));
    layer0_outputs(7817) <= (inputs(189)) or (inputs(219));
    layer0_outputs(7818) <= '0';
    layer0_outputs(7819) <= not((inputs(97)) and (inputs(120)));
    layer0_outputs(7820) <= not((inputs(155)) xor (inputs(238)));
    layer0_outputs(7821) <= not(inputs(7));
    layer0_outputs(7822) <= not((inputs(201)) or (inputs(41)));
    layer0_outputs(7823) <= not((inputs(223)) or (inputs(214)));
    layer0_outputs(7824) <= inputs(174);
    layer0_outputs(7825) <= (inputs(9)) and not (inputs(87));
    layer0_outputs(7826) <= not((inputs(99)) or (inputs(47)));
    layer0_outputs(7827) <= not(inputs(165));
    layer0_outputs(7828) <= '1';
    layer0_outputs(7829) <= not((inputs(43)) xor (inputs(30)));
    layer0_outputs(7830) <= not((inputs(235)) or (inputs(147)));
    layer0_outputs(7831) <= inputs(186);
    layer0_outputs(7832) <= not((inputs(108)) xor (inputs(28)));
    layer0_outputs(7833) <= not((inputs(221)) xor (inputs(15)));
    layer0_outputs(7834) <= not(inputs(214));
    layer0_outputs(7835) <= (inputs(122)) and not (inputs(11));
    layer0_outputs(7836) <= inputs(253);
    layer0_outputs(7837) <= not((inputs(203)) and (inputs(201)));
    layer0_outputs(7838) <= not(inputs(157)) or (inputs(132));
    layer0_outputs(7839) <= inputs(82);
    layer0_outputs(7840) <= not(inputs(213));
    layer0_outputs(7841) <= inputs(141);
    layer0_outputs(7842) <= not(inputs(94));
    layer0_outputs(7843) <= not(inputs(68));
    layer0_outputs(7844) <= not((inputs(235)) or (inputs(134)));
    layer0_outputs(7845) <= (inputs(197)) and not (inputs(41));
    layer0_outputs(7846) <= (inputs(65)) or (inputs(159));
    layer0_outputs(7847) <= not(inputs(88));
    layer0_outputs(7848) <= inputs(83);
    layer0_outputs(7849) <= not((inputs(36)) xor (inputs(187)));
    layer0_outputs(7850) <= not(inputs(230));
    layer0_outputs(7851) <= (inputs(140)) and not (inputs(98));
    layer0_outputs(7852) <= inputs(153);
    layer0_outputs(7853) <= (inputs(133)) and not (inputs(172));
    layer0_outputs(7854) <= inputs(40);
    layer0_outputs(7855) <= (inputs(170)) xor (inputs(234));
    layer0_outputs(7856) <= not(inputs(153));
    layer0_outputs(7857) <= (inputs(224)) or (inputs(17));
    layer0_outputs(7858) <= (inputs(221)) and not (inputs(143));
    layer0_outputs(7859) <= not(inputs(134)) or (inputs(222));
    layer0_outputs(7860) <= inputs(234);
    layer0_outputs(7861) <= not(inputs(230));
    layer0_outputs(7862) <= (inputs(225)) and not (inputs(193));
    layer0_outputs(7863) <= not(inputs(135)) or (inputs(176));
    layer0_outputs(7864) <= not((inputs(197)) or (inputs(141)));
    layer0_outputs(7865) <= not(inputs(132)) or (inputs(242));
    layer0_outputs(7866) <= (inputs(208)) xor (inputs(126));
    layer0_outputs(7867) <= (inputs(150)) and not (inputs(245));
    layer0_outputs(7868) <= not(inputs(55)) or (inputs(4));
    layer0_outputs(7869) <= not((inputs(58)) or (inputs(24)));
    layer0_outputs(7870) <= not(inputs(4));
    layer0_outputs(7871) <= not(inputs(215)) or (inputs(35));
    layer0_outputs(7872) <= inputs(32);
    layer0_outputs(7873) <= (inputs(173)) or (inputs(250));
    layer0_outputs(7874) <= inputs(165);
    layer0_outputs(7875) <= not(inputs(155)) or (inputs(105));
    layer0_outputs(7876) <= (inputs(185)) and not (inputs(56));
    layer0_outputs(7877) <= inputs(24);
    layer0_outputs(7878) <= (inputs(32)) or (inputs(123));
    layer0_outputs(7879) <= not(inputs(108));
    layer0_outputs(7880) <= not(inputs(237));
    layer0_outputs(7881) <= (inputs(119)) and not (inputs(207));
    layer0_outputs(7882) <= (inputs(143)) xor (inputs(191));
    layer0_outputs(7883) <= (inputs(153)) and not (inputs(105));
    layer0_outputs(7884) <= inputs(87);
    layer0_outputs(7885) <= (inputs(255)) or (inputs(197));
    layer0_outputs(7886) <= (inputs(156)) and not (inputs(0));
    layer0_outputs(7887) <= not((inputs(72)) or (inputs(131)));
    layer0_outputs(7888) <= not((inputs(169)) or (inputs(177)));
    layer0_outputs(7889) <= inputs(168);
    layer0_outputs(7890) <= inputs(111);
    layer0_outputs(7891) <= (inputs(53)) and not (inputs(246));
    layer0_outputs(7892) <= inputs(91);
    layer0_outputs(7893) <= not(inputs(105));
    layer0_outputs(7894) <= not((inputs(234)) or (inputs(161)));
    layer0_outputs(7895) <= (inputs(208)) and (inputs(250));
    layer0_outputs(7896) <= (inputs(200)) and not (inputs(106));
    layer0_outputs(7897) <= not(inputs(229)) or (inputs(99));
    layer0_outputs(7898) <= (inputs(239)) or (inputs(66));
    layer0_outputs(7899) <= not((inputs(65)) or (inputs(152)));
    layer0_outputs(7900) <= not((inputs(30)) or (inputs(154)));
    layer0_outputs(7901) <= not(inputs(148));
    layer0_outputs(7902) <= inputs(23);
    layer0_outputs(7903) <= (inputs(21)) and not (inputs(126));
    layer0_outputs(7904) <= '0';
    layer0_outputs(7905) <= (inputs(224)) or (inputs(201));
    layer0_outputs(7906) <= inputs(212);
    layer0_outputs(7907) <= not(inputs(115)) or (inputs(204));
    layer0_outputs(7908) <= (inputs(89)) and not (inputs(224));
    layer0_outputs(7909) <= not((inputs(215)) or (inputs(119)));
    layer0_outputs(7910) <= '0';
    layer0_outputs(7911) <= '0';
    layer0_outputs(7912) <= inputs(106);
    layer0_outputs(7913) <= (inputs(102)) xor (inputs(10));
    layer0_outputs(7914) <= not((inputs(157)) and (inputs(37)));
    layer0_outputs(7915) <= (inputs(117)) and (inputs(13));
    layer0_outputs(7916) <= '0';
    layer0_outputs(7917) <= not((inputs(161)) or (inputs(32)));
    layer0_outputs(7918) <= not(inputs(126));
    layer0_outputs(7919) <= (inputs(135)) or (inputs(47));
    layer0_outputs(7920) <= not((inputs(164)) or (inputs(162)));
    layer0_outputs(7921) <= not((inputs(24)) or (inputs(64)));
    layer0_outputs(7922) <= not((inputs(164)) or (inputs(81)));
    layer0_outputs(7923) <= (inputs(182)) or (inputs(96));
    layer0_outputs(7924) <= not(inputs(239)) or (inputs(81));
    layer0_outputs(7925) <= not(inputs(65)) or (inputs(21));
    layer0_outputs(7926) <= not(inputs(244)) or (inputs(111));
    layer0_outputs(7927) <= not(inputs(236)) or (inputs(140));
    layer0_outputs(7928) <= (inputs(230)) or (inputs(94));
    layer0_outputs(7929) <= (inputs(101)) and not (inputs(219));
    layer0_outputs(7930) <= (inputs(151)) and not (inputs(82));
    layer0_outputs(7931) <= (inputs(120)) xor (inputs(219));
    layer0_outputs(7932) <= inputs(184);
    layer0_outputs(7933) <= (inputs(248)) and not (inputs(50));
    layer0_outputs(7934) <= not((inputs(141)) and (inputs(210)));
    layer0_outputs(7935) <= (inputs(182)) and not (inputs(11));
    layer0_outputs(7936) <= '1';
    layer0_outputs(7937) <= not((inputs(86)) or (inputs(87)));
    layer0_outputs(7938) <= inputs(233);
    layer0_outputs(7939) <= not(inputs(106));
    layer0_outputs(7940) <= not(inputs(121));
    layer0_outputs(7941) <= (inputs(16)) or (inputs(97));
    layer0_outputs(7942) <= (inputs(233)) and not (inputs(116));
    layer0_outputs(7943) <= (inputs(142)) and not (inputs(237));
    layer0_outputs(7944) <= inputs(144);
    layer0_outputs(7945) <= inputs(148);
    layer0_outputs(7946) <= inputs(97);
    layer0_outputs(7947) <= inputs(131);
    layer0_outputs(7948) <= not(inputs(194)) or (inputs(45));
    layer0_outputs(7949) <= not(inputs(217));
    layer0_outputs(7950) <= (inputs(224)) or (inputs(168));
    layer0_outputs(7951) <= '0';
    layer0_outputs(7952) <= not(inputs(52));
    layer0_outputs(7953) <= (inputs(115)) xor (inputs(52));
    layer0_outputs(7954) <= not(inputs(58)) or (inputs(214));
    layer0_outputs(7955) <= not((inputs(108)) or (inputs(37)));
    layer0_outputs(7956) <= inputs(216);
    layer0_outputs(7957) <= not((inputs(199)) xor (inputs(247)));
    layer0_outputs(7958) <= (inputs(212)) or (inputs(23));
    layer0_outputs(7959) <= not(inputs(103)) or (inputs(125));
    layer0_outputs(7960) <= not((inputs(49)) or (inputs(249)));
    layer0_outputs(7961) <= (inputs(236)) or (inputs(18));
    layer0_outputs(7962) <= not((inputs(195)) or (inputs(178)));
    layer0_outputs(7963) <= inputs(254);
    layer0_outputs(7964) <= inputs(44);
    layer0_outputs(7965) <= not(inputs(208)) or (inputs(190));
    layer0_outputs(7966) <= (inputs(139)) xor (inputs(252));
    layer0_outputs(7967) <= (inputs(35)) or (inputs(195));
    layer0_outputs(7968) <= not((inputs(160)) or (inputs(152)));
    layer0_outputs(7969) <= (inputs(147)) or (inputs(130));
    layer0_outputs(7970) <= not(inputs(218)) or (inputs(231));
    layer0_outputs(7971) <= inputs(141);
    layer0_outputs(7972) <= not((inputs(115)) xor (inputs(128)));
    layer0_outputs(7973) <= not((inputs(87)) or (inputs(135)));
    layer0_outputs(7974) <= (inputs(210)) or (inputs(114));
    layer0_outputs(7975) <= (inputs(165)) and not (inputs(207));
    layer0_outputs(7976) <= (inputs(142)) or (inputs(2));
    layer0_outputs(7977) <= (inputs(228)) xor (inputs(254));
    layer0_outputs(7978) <= (inputs(65)) and not (inputs(45));
    layer0_outputs(7979) <= (inputs(94)) or (inputs(149));
    layer0_outputs(7980) <= not((inputs(166)) or (inputs(44)));
    layer0_outputs(7981) <= (inputs(107)) and not (inputs(81));
    layer0_outputs(7982) <= '0';
    layer0_outputs(7983) <= (inputs(209)) and not (inputs(1));
    layer0_outputs(7984) <= not((inputs(88)) xor (inputs(118)));
    layer0_outputs(7985) <= not((inputs(206)) xor (inputs(97)));
    layer0_outputs(7986) <= '1';
    layer0_outputs(7987) <= (inputs(75)) or (inputs(107));
    layer0_outputs(7988) <= '1';
    layer0_outputs(7989) <= not(inputs(233));
    layer0_outputs(7990) <= inputs(119);
    layer0_outputs(7991) <= (inputs(5)) and not (inputs(186));
    layer0_outputs(7992) <= not((inputs(202)) and (inputs(75)));
    layer0_outputs(7993) <= not(inputs(183)) or (inputs(48));
    layer0_outputs(7994) <= not(inputs(105)) or (inputs(140));
    layer0_outputs(7995) <= not(inputs(198));
    layer0_outputs(7996) <= '0';
    layer0_outputs(7997) <= not(inputs(39)) or (inputs(178));
    layer0_outputs(7998) <= (inputs(100)) xor (inputs(3));
    layer0_outputs(7999) <= not(inputs(82));
    layer0_outputs(8000) <= (inputs(182)) and not (inputs(72));
    layer0_outputs(8001) <= not(inputs(109));
    layer0_outputs(8002) <= not(inputs(251));
    layer0_outputs(8003) <= not(inputs(3)) or (inputs(175));
    layer0_outputs(8004) <= inputs(10);
    layer0_outputs(8005) <= (inputs(205)) xor (inputs(125));
    layer0_outputs(8006) <= not(inputs(206));
    layer0_outputs(8007) <= inputs(151);
    layer0_outputs(8008) <= (inputs(140)) and not (inputs(163));
    layer0_outputs(8009) <= (inputs(111)) xor (inputs(140));
    layer0_outputs(8010) <= not(inputs(7));
    layer0_outputs(8011) <= not((inputs(63)) or (inputs(10)));
    layer0_outputs(8012) <= inputs(231);
    layer0_outputs(8013) <= not(inputs(164));
    layer0_outputs(8014) <= (inputs(146)) or (inputs(81));
    layer0_outputs(8015) <= (inputs(147)) or (inputs(2));
    layer0_outputs(8016) <= not((inputs(223)) or (inputs(39)));
    layer0_outputs(8017) <= not(inputs(19));
    layer0_outputs(8018) <= not(inputs(54)) or (inputs(31));
    layer0_outputs(8019) <= (inputs(183)) and not (inputs(176));
    layer0_outputs(8020) <= not(inputs(192)) or (inputs(221));
    layer0_outputs(8021) <= not((inputs(20)) or (inputs(230)));
    layer0_outputs(8022) <= inputs(80);
    layer0_outputs(8023) <= (inputs(252)) and not (inputs(224));
    layer0_outputs(8024) <= inputs(229);
    layer0_outputs(8025) <= inputs(112);
    layer0_outputs(8026) <= inputs(163);
    layer0_outputs(8027) <= inputs(237);
    layer0_outputs(8028) <= not((inputs(128)) xor (inputs(70)));
    layer0_outputs(8029) <= '0';
    layer0_outputs(8030) <= '0';
    layer0_outputs(8031) <= not(inputs(229));
    layer0_outputs(8032) <= '0';
    layer0_outputs(8033) <= (inputs(135)) or (inputs(49));
    layer0_outputs(8034) <= (inputs(176)) or (inputs(246));
    layer0_outputs(8035) <= not(inputs(137));
    layer0_outputs(8036) <= not(inputs(53)) or (inputs(154));
    layer0_outputs(8037) <= inputs(152);
    layer0_outputs(8038) <= (inputs(62)) xor (inputs(24));
    layer0_outputs(8039) <= (inputs(1)) or (inputs(226));
    layer0_outputs(8040) <= inputs(193);
    layer0_outputs(8041) <= not(inputs(250));
    layer0_outputs(8042) <= not(inputs(199)) or (inputs(28));
    layer0_outputs(8043) <= inputs(15);
    layer0_outputs(8044) <= not(inputs(108)) or (inputs(34));
    layer0_outputs(8045) <= inputs(194);
    layer0_outputs(8046) <= inputs(95);
    layer0_outputs(8047) <= (inputs(23)) xor (inputs(0));
    layer0_outputs(8048) <= (inputs(120)) and (inputs(242));
    layer0_outputs(8049) <= not(inputs(19)) or (inputs(28));
    layer0_outputs(8050) <= inputs(69);
    layer0_outputs(8051) <= inputs(171);
    layer0_outputs(8052) <= (inputs(54)) and not (inputs(91));
    layer0_outputs(8053) <= not(inputs(43));
    layer0_outputs(8054) <= (inputs(249)) and not (inputs(63));
    layer0_outputs(8055) <= not((inputs(6)) or (inputs(27)));
    layer0_outputs(8056) <= not(inputs(118)) or (inputs(65));
    layer0_outputs(8057) <= not((inputs(57)) or (inputs(16)));
    layer0_outputs(8058) <= not((inputs(82)) or (inputs(22)));
    layer0_outputs(8059) <= not((inputs(64)) or (inputs(50)));
    layer0_outputs(8060) <= not((inputs(124)) or (inputs(129)));
    layer0_outputs(8061) <= not((inputs(253)) or (inputs(206)));
    layer0_outputs(8062) <= inputs(171);
    layer0_outputs(8063) <= not(inputs(246));
    layer0_outputs(8064) <= (inputs(23)) and not (inputs(29));
    layer0_outputs(8065) <= not(inputs(220));
    layer0_outputs(8066) <= '1';
    layer0_outputs(8067) <= not(inputs(90));
    layer0_outputs(8068) <= inputs(113);
    layer0_outputs(8069) <= not(inputs(197));
    layer0_outputs(8070) <= '1';
    layer0_outputs(8071) <= not(inputs(236)) or (inputs(110));
    layer0_outputs(8072) <= not(inputs(163)) or (inputs(24));
    layer0_outputs(8073) <= inputs(221);
    layer0_outputs(8074) <= not(inputs(169)) or (inputs(105));
    layer0_outputs(8075) <= not((inputs(245)) and (inputs(217)));
    layer0_outputs(8076) <= not(inputs(165));
    layer0_outputs(8077) <= not(inputs(83)) or (inputs(194));
    layer0_outputs(8078) <= (inputs(236)) or (inputs(69));
    layer0_outputs(8079) <= (inputs(147)) and not (inputs(104));
    layer0_outputs(8080) <= (inputs(95)) and (inputs(254));
    layer0_outputs(8081) <= not(inputs(131));
    layer0_outputs(8082) <= (inputs(47)) or (inputs(143));
    layer0_outputs(8083) <= inputs(175);
    layer0_outputs(8084) <= not(inputs(54)) or (inputs(129));
    layer0_outputs(8085) <= (inputs(73)) and not (inputs(2));
    layer0_outputs(8086) <= not(inputs(90));
    layer0_outputs(8087) <= not(inputs(84));
    layer0_outputs(8088) <= not(inputs(146));
    layer0_outputs(8089) <= (inputs(47)) and (inputs(227));
    layer0_outputs(8090) <= not((inputs(216)) or (inputs(137)));
    layer0_outputs(8091) <= inputs(94);
    layer0_outputs(8092) <= inputs(202);
    layer0_outputs(8093) <= inputs(165);
    layer0_outputs(8094) <= not(inputs(121)) or (inputs(207));
    layer0_outputs(8095) <= not(inputs(167)) or (inputs(145));
    layer0_outputs(8096) <= inputs(8);
    layer0_outputs(8097) <= (inputs(42)) and not (inputs(236));
    layer0_outputs(8098) <= not(inputs(148));
    layer0_outputs(8099) <= not(inputs(246));
    layer0_outputs(8100) <= not(inputs(53)) or (inputs(225));
    layer0_outputs(8101) <= not(inputs(37));
    layer0_outputs(8102) <= not(inputs(235)) or (inputs(138));
    layer0_outputs(8103) <= (inputs(76)) or (inputs(37));
    layer0_outputs(8104) <= (inputs(54)) or (inputs(165));
    layer0_outputs(8105) <= (inputs(158)) or (inputs(12));
    layer0_outputs(8106) <= not(inputs(133)) or (inputs(18));
    layer0_outputs(8107) <= not(inputs(38)) or (inputs(116));
    layer0_outputs(8108) <= not(inputs(144));
    layer0_outputs(8109) <= (inputs(30)) and not (inputs(29));
    layer0_outputs(8110) <= '0';
    layer0_outputs(8111) <= not((inputs(107)) xor (inputs(19)));
    layer0_outputs(8112) <= inputs(82);
    layer0_outputs(8113) <= not((inputs(207)) and (inputs(245)));
    layer0_outputs(8114) <= not(inputs(182)) or (inputs(78));
    layer0_outputs(8115) <= (inputs(20)) and not (inputs(109));
    layer0_outputs(8116) <= (inputs(168)) or (inputs(23));
    layer0_outputs(8117) <= not(inputs(65)) or (inputs(1));
    layer0_outputs(8118) <= not(inputs(100)) or (inputs(57));
    layer0_outputs(8119) <= not((inputs(18)) and (inputs(47)));
    layer0_outputs(8120) <= (inputs(166)) or (inputs(191));
    layer0_outputs(8121) <= inputs(94);
    layer0_outputs(8122) <= (inputs(205)) and not (inputs(167));
    layer0_outputs(8123) <= not((inputs(40)) xor (inputs(31)));
    layer0_outputs(8124) <= not(inputs(55)) or (inputs(45));
    layer0_outputs(8125) <= '0';
    layer0_outputs(8126) <= not(inputs(149)) or (inputs(222));
    layer0_outputs(8127) <= not(inputs(200));
    layer0_outputs(8128) <= inputs(253);
    layer0_outputs(8129) <= not((inputs(246)) or (inputs(176)));
    layer0_outputs(8130) <= not(inputs(183)) or (inputs(48));
    layer0_outputs(8131) <= not(inputs(115)) or (inputs(62));
    layer0_outputs(8132) <= '1';
    layer0_outputs(8133) <= (inputs(6)) xor (inputs(31));
    layer0_outputs(8134) <= inputs(192);
    layer0_outputs(8135) <= not((inputs(181)) or (inputs(208)));
    layer0_outputs(8136) <= (inputs(200)) or (inputs(163));
    layer0_outputs(8137) <= '0';
    layer0_outputs(8138) <= not(inputs(202));
    layer0_outputs(8139) <= (inputs(245)) and not (inputs(110));
    layer0_outputs(8140) <= (inputs(16)) xor (inputs(108));
    layer0_outputs(8141) <= not(inputs(78));
    layer0_outputs(8142) <= not(inputs(89));
    layer0_outputs(8143) <= not(inputs(10));
    layer0_outputs(8144) <= (inputs(100)) and not (inputs(219));
    layer0_outputs(8145) <= not(inputs(96)) or (inputs(208));
    layer0_outputs(8146) <= not((inputs(207)) xor (inputs(209)));
    layer0_outputs(8147) <= not((inputs(88)) or (inputs(60)));
    layer0_outputs(8148) <= not((inputs(225)) or (inputs(110)));
    layer0_outputs(8149) <= not((inputs(62)) or (inputs(151)));
    layer0_outputs(8150) <= not((inputs(221)) or (inputs(218)));
    layer0_outputs(8151) <= (inputs(156)) and (inputs(169));
    layer0_outputs(8152) <= (inputs(95)) xor (inputs(75));
    layer0_outputs(8153) <= not((inputs(176)) xor (inputs(170)));
    layer0_outputs(8154) <= not(inputs(205)) or (inputs(79));
    layer0_outputs(8155) <= (inputs(131)) or (inputs(239));
    layer0_outputs(8156) <= not((inputs(73)) xor (inputs(24)));
    layer0_outputs(8157) <= not(inputs(209));
    layer0_outputs(8158) <= (inputs(229)) and not (inputs(78));
    layer0_outputs(8159) <= (inputs(32)) or (inputs(45));
    layer0_outputs(8160) <= not(inputs(117));
    layer0_outputs(8161) <= not(inputs(231));
    layer0_outputs(8162) <= inputs(75);
    layer0_outputs(8163) <= not(inputs(178));
    layer0_outputs(8164) <= not((inputs(182)) and (inputs(177)));
    layer0_outputs(8165) <= (inputs(46)) xor (inputs(14));
    layer0_outputs(8166) <= inputs(237);
    layer0_outputs(8167) <= '0';
    layer0_outputs(8168) <= (inputs(128)) and not (inputs(61));
    layer0_outputs(8169) <= (inputs(83)) or (inputs(154));
    layer0_outputs(8170) <= not((inputs(192)) and (inputs(212)));
    layer0_outputs(8171) <= inputs(162);
    layer0_outputs(8172) <= '1';
    layer0_outputs(8173) <= (inputs(136)) and not (inputs(51));
    layer0_outputs(8174) <= (inputs(75)) and not (inputs(117));
    layer0_outputs(8175) <= inputs(26);
    layer0_outputs(8176) <= not(inputs(74)) or (inputs(223));
    layer0_outputs(8177) <= (inputs(120)) or (inputs(236));
    layer0_outputs(8178) <= (inputs(248)) and (inputs(114));
    layer0_outputs(8179) <= inputs(55);
    layer0_outputs(8180) <= '1';
    layer0_outputs(8181) <= not(inputs(75)) or (inputs(252));
    layer0_outputs(8182) <= (inputs(158)) and (inputs(102));
    layer0_outputs(8183) <= (inputs(34)) and (inputs(47));
    layer0_outputs(8184) <= inputs(170);
    layer0_outputs(8185) <= inputs(113);
    layer0_outputs(8186) <= not(inputs(112));
    layer0_outputs(8187) <= (inputs(197)) and not (inputs(140));
    layer0_outputs(8188) <= (inputs(127)) and not (inputs(49));
    layer0_outputs(8189) <= '0';
    layer0_outputs(8190) <= not((inputs(4)) or (inputs(177)));
    layer0_outputs(8191) <= not(inputs(63));
    layer0_outputs(8192) <= (inputs(239)) xor (inputs(84));
    layer0_outputs(8193) <= (inputs(34)) and (inputs(219));
    layer0_outputs(8194) <= not(inputs(34));
    layer0_outputs(8195) <= inputs(158);
    layer0_outputs(8196) <= inputs(40);
    layer0_outputs(8197) <= (inputs(166)) or (inputs(252));
    layer0_outputs(8198) <= not(inputs(113));
    layer0_outputs(8199) <= not((inputs(173)) or (inputs(42)));
    layer0_outputs(8200) <= not(inputs(81)) or (inputs(196));
    layer0_outputs(8201) <= not(inputs(104));
    layer0_outputs(8202) <= (inputs(168)) and not (inputs(251));
    layer0_outputs(8203) <= not(inputs(153));
    layer0_outputs(8204) <= (inputs(108)) and (inputs(153));
    layer0_outputs(8205) <= not((inputs(33)) or (inputs(200)));
    layer0_outputs(8206) <= (inputs(130)) xor (inputs(162));
    layer0_outputs(8207) <= not((inputs(135)) or (inputs(22)));
    layer0_outputs(8208) <= inputs(133);
    layer0_outputs(8209) <= (inputs(157)) and not (inputs(231));
    layer0_outputs(8210) <= not(inputs(105));
    layer0_outputs(8211) <= not(inputs(164));
    layer0_outputs(8212) <= not((inputs(155)) xor (inputs(8)));
    layer0_outputs(8213) <= inputs(210);
    layer0_outputs(8214) <= inputs(126);
    layer0_outputs(8215) <= not(inputs(35));
    layer0_outputs(8216) <= (inputs(148)) and not (inputs(160));
    layer0_outputs(8217) <= not((inputs(221)) or (inputs(48)));
    layer0_outputs(8218) <= (inputs(171)) and not (inputs(211));
    layer0_outputs(8219) <= not((inputs(191)) xor (inputs(70)));
    layer0_outputs(8220) <= not(inputs(56)) or (inputs(233));
    layer0_outputs(8221) <= not(inputs(160)) or (inputs(112));
    layer0_outputs(8222) <= (inputs(223)) xor (inputs(28));
    layer0_outputs(8223) <= (inputs(222)) xor (inputs(221));
    layer0_outputs(8224) <= not(inputs(122));
    layer0_outputs(8225) <= not(inputs(25));
    layer0_outputs(8226) <= inputs(167);
    layer0_outputs(8227) <= not((inputs(221)) or (inputs(205)));
    layer0_outputs(8228) <= (inputs(216)) xor (inputs(176));
    layer0_outputs(8229) <= not(inputs(217));
    layer0_outputs(8230) <= inputs(79);
    layer0_outputs(8231) <= (inputs(106)) and not (inputs(17));
    layer0_outputs(8232) <= not(inputs(199)) or (inputs(108));
    layer0_outputs(8233) <= inputs(207);
    layer0_outputs(8234) <= not(inputs(38)) or (inputs(73));
    layer0_outputs(8235) <= not((inputs(199)) or (inputs(237)));
    layer0_outputs(8236) <= inputs(75);
    layer0_outputs(8237) <= (inputs(190)) or (inputs(174));
    layer0_outputs(8238) <= (inputs(104)) or (inputs(2));
    layer0_outputs(8239) <= not(inputs(198));
    layer0_outputs(8240) <= inputs(94);
    layer0_outputs(8241) <= (inputs(2)) or (inputs(38));
    layer0_outputs(8242) <= not(inputs(59)) or (inputs(254));
    layer0_outputs(8243) <= (inputs(79)) and (inputs(80));
    layer0_outputs(8244) <= not(inputs(123)) or (inputs(196));
    layer0_outputs(8245) <= (inputs(30)) and (inputs(254));
    layer0_outputs(8246) <= not(inputs(211));
    layer0_outputs(8247) <= (inputs(124)) and not (inputs(14));
    layer0_outputs(8248) <= not(inputs(146));
    layer0_outputs(8249) <= not(inputs(210)) or (inputs(99));
    layer0_outputs(8250) <= (inputs(9)) xor (inputs(116));
    layer0_outputs(8251) <= (inputs(229)) or (inputs(102));
    layer0_outputs(8252) <= not((inputs(206)) or (inputs(32)));
    layer0_outputs(8253) <= (inputs(118)) or (inputs(175));
    layer0_outputs(8254) <= (inputs(66)) and not (inputs(190));
    layer0_outputs(8255) <= not((inputs(179)) xor (inputs(127)));
    layer0_outputs(8256) <= '0';
    layer0_outputs(8257) <= '1';
    layer0_outputs(8258) <= inputs(86);
    layer0_outputs(8259) <= not(inputs(220)) or (inputs(12));
    layer0_outputs(8260) <= (inputs(103)) and not (inputs(237));
    layer0_outputs(8261) <= not((inputs(39)) or (inputs(205)));
    layer0_outputs(8262) <= not(inputs(96));
    layer0_outputs(8263) <= not((inputs(154)) xor (inputs(203)));
    layer0_outputs(8264) <= not((inputs(188)) or (inputs(57)));
    layer0_outputs(8265) <= not((inputs(237)) or (inputs(188)));
    layer0_outputs(8266) <= not(inputs(37)) or (inputs(84));
    layer0_outputs(8267) <= inputs(40);
    layer0_outputs(8268) <= not((inputs(196)) or (inputs(162)));
    layer0_outputs(8269) <= (inputs(180)) and not (inputs(4));
    layer0_outputs(8270) <= (inputs(95)) and not (inputs(16));
    layer0_outputs(8271) <= '0';
    layer0_outputs(8272) <= (inputs(0)) and not (inputs(172));
    layer0_outputs(8273) <= not(inputs(147));
    layer0_outputs(8274) <= '0';
    layer0_outputs(8275) <= not((inputs(92)) or (inputs(115)));
    layer0_outputs(8276) <= not(inputs(183)) or (inputs(113));
    layer0_outputs(8277) <= '1';
    layer0_outputs(8278) <= not(inputs(119));
    layer0_outputs(8279) <= not(inputs(239)) or (inputs(233));
    layer0_outputs(8280) <= inputs(238);
    layer0_outputs(8281) <= (inputs(159)) xor (inputs(117));
    layer0_outputs(8282) <= not(inputs(62));
    layer0_outputs(8283) <= not((inputs(236)) and (inputs(214)));
    layer0_outputs(8284) <= not((inputs(130)) or (inputs(162)));
    layer0_outputs(8285) <= '1';
    layer0_outputs(8286) <= not(inputs(102)) or (inputs(16));
    layer0_outputs(8287) <= not((inputs(17)) xor (inputs(140)));
    layer0_outputs(8288) <= not(inputs(50));
    layer0_outputs(8289) <= (inputs(27)) xor (inputs(59));
    layer0_outputs(8290) <= (inputs(89)) xor (inputs(55));
    layer0_outputs(8291) <= '1';
    layer0_outputs(8292) <= (inputs(238)) and not (inputs(39));
    layer0_outputs(8293) <= not((inputs(174)) or (inputs(29)));
    layer0_outputs(8294) <= not(inputs(83)) or (inputs(162));
    layer0_outputs(8295) <= not(inputs(57));
    layer0_outputs(8296) <= not((inputs(170)) and (inputs(209)));
    layer0_outputs(8297) <= (inputs(164)) xor (inputs(203));
    layer0_outputs(8298) <= (inputs(166)) xor (inputs(50));
    layer0_outputs(8299) <= inputs(191);
    layer0_outputs(8300) <= (inputs(114)) and (inputs(138));
    layer0_outputs(8301) <= inputs(144);
    layer0_outputs(8302) <= not(inputs(75));
    layer0_outputs(8303) <= (inputs(168)) and not (inputs(77));
    layer0_outputs(8304) <= not(inputs(178));
    layer0_outputs(8305) <= '1';
    layer0_outputs(8306) <= (inputs(89)) xor (inputs(84));
    layer0_outputs(8307) <= not((inputs(39)) xor (inputs(143)));
    layer0_outputs(8308) <= inputs(76);
    layer0_outputs(8309) <= inputs(116);
    layer0_outputs(8310) <= (inputs(212)) or (inputs(63));
    layer0_outputs(8311) <= inputs(111);
    layer0_outputs(8312) <= inputs(201);
    layer0_outputs(8313) <= not(inputs(188)) or (inputs(19));
    layer0_outputs(8314) <= not(inputs(20));
    layer0_outputs(8315) <= not(inputs(181)) or (inputs(117));
    layer0_outputs(8316) <= not(inputs(250)) or (inputs(20));
    layer0_outputs(8317) <= not(inputs(177));
    layer0_outputs(8318) <= (inputs(136)) xor (inputs(89));
    layer0_outputs(8319) <= (inputs(146)) and (inputs(102));
    layer0_outputs(8320) <= inputs(118);
    layer0_outputs(8321) <= not((inputs(241)) or (inputs(110)));
    layer0_outputs(8322) <= inputs(26);
    layer0_outputs(8323) <= not((inputs(69)) xor (inputs(2)));
    layer0_outputs(8324) <= '1';
    layer0_outputs(8325) <= (inputs(123)) or (inputs(135));
    layer0_outputs(8326) <= not((inputs(176)) or (inputs(116)));
    layer0_outputs(8327) <= not(inputs(67));
    layer0_outputs(8328) <= not(inputs(113)) or (inputs(87));
    layer0_outputs(8329) <= not(inputs(204));
    layer0_outputs(8330) <= (inputs(149)) or (inputs(153));
    layer0_outputs(8331) <= inputs(129);
    layer0_outputs(8332) <= not(inputs(68)) or (inputs(33));
    layer0_outputs(8333) <= inputs(154);
    layer0_outputs(8334) <= inputs(147);
    layer0_outputs(8335) <= (inputs(141)) and not (inputs(18));
    layer0_outputs(8336) <= not((inputs(93)) or (inputs(226)));
    layer0_outputs(8337) <= not((inputs(159)) xor (inputs(216)));
    layer0_outputs(8338) <= (inputs(154)) or (inputs(219));
    layer0_outputs(8339) <= inputs(151);
    layer0_outputs(8340) <= not(inputs(10));
    layer0_outputs(8341) <= not((inputs(180)) or (inputs(6)));
    layer0_outputs(8342) <= not(inputs(40));
    layer0_outputs(8343) <= not(inputs(228)) or (inputs(30));
    layer0_outputs(8344) <= (inputs(65)) and not (inputs(202));
    layer0_outputs(8345) <= not(inputs(106));
    layer0_outputs(8346) <= inputs(232);
    layer0_outputs(8347) <= not(inputs(98));
    layer0_outputs(8348) <= inputs(120);
    layer0_outputs(8349) <= inputs(162);
    layer0_outputs(8350) <= '0';
    layer0_outputs(8351) <= '1';
    layer0_outputs(8352) <= not((inputs(203)) or (inputs(129)));
    layer0_outputs(8353) <= (inputs(178)) or (inputs(109));
    layer0_outputs(8354) <= not(inputs(43)) or (inputs(190));
    layer0_outputs(8355) <= inputs(166);
    layer0_outputs(8356) <= (inputs(212)) and not (inputs(36));
    layer0_outputs(8357) <= (inputs(240)) xor (inputs(237));
    layer0_outputs(8358) <= inputs(25);
    layer0_outputs(8359) <= inputs(124);
    layer0_outputs(8360) <= not(inputs(4));
    layer0_outputs(8361) <= (inputs(116)) and not (inputs(226));
    layer0_outputs(8362) <= (inputs(108)) xor (inputs(169));
    layer0_outputs(8363) <= inputs(82);
    layer0_outputs(8364) <= not(inputs(47)) or (inputs(109));
    layer0_outputs(8365) <= not(inputs(247));
    layer0_outputs(8366) <= inputs(102);
    layer0_outputs(8367) <= (inputs(91)) and (inputs(251));
    layer0_outputs(8368) <= not((inputs(130)) or (inputs(112)));
    layer0_outputs(8369) <= not(inputs(207)) or (inputs(226));
    layer0_outputs(8370) <= not(inputs(187));
    layer0_outputs(8371) <= inputs(160);
    layer0_outputs(8372) <= not(inputs(124));
    layer0_outputs(8373) <= inputs(201);
    layer0_outputs(8374) <= not((inputs(58)) or (inputs(16)));
    layer0_outputs(8375) <= inputs(138);
    layer0_outputs(8376) <= inputs(237);
    layer0_outputs(8377) <= (inputs(87)) and not (inputs(233));
    layer0_outputs(8378) <= (inputs(33)) or (inputs(57));
    layer0_outputs(8379) <= (inputs(220)) or (inputs(127));
    layer0_outputs(8380) <= (inputs(34)) and (inputs(93));
    layer0_outputs(8381) <= not((inputs(124)) or (inputs(190)));
    layer0_outputs(8382) <= not(inputs(148)) or (inputs(191));
    layer0_outputs(8383) <= (inputs(26)) and not (inputs(151));
    layer0_outputs(8384) <= inputs(116);
    layer0_outputs(8385) <= not((inputs(0)) xor (inputs(211)));
    layer0_outputs(8386) <= not(inputs(253));
    layer0_outputs(8387) <= not(inputs(97));
    layer0_outputs(8388) <= (inputs(154)) and (inputs(87));
    layer0_outputs(8389) <= not(inputs(2)) or (inputs(232));
    layer0_outputs(8390) <= not((inputs(160)) or (inputs(213)));
    layer0_outputs(8391) <= (inputs(64)) or (inputs(205));
    layer0_outputs(8392) <= inputs(104);
    layer0_outputs(8393) <= inputs(59);
    layer0_outputs(8394) <= not((inputs(19)) xor (inputs(50)));
    layer0_outputs(8395) <= (inputs(224)) and not (inputs(103));
    layer0_outputs(8396) <= not(inputs(35)) or (inputs(139));
    layer0_outputs(8397) <= not((inputs(16)) xor (inputs(225)));
    layer0_outputs(8398) <= (inputs(13)) xor (inputs(127));
    layer0_outputs(8399) <= (inputs(221)) and not (inputs(15));
    layer0_outputs(8400) <= '0';
    layer0_outputs(8401) <= not((inputs(193)) or (inputs(176)));
    layer0_outputs(8402) <= not(inputs(155)) or (inputs(188));
    layer0_outputs(8403) <= inputs(89);
    layer0_outputs(8404) <= inputs(118);
    layer0_outputs(8405) <= not(inputs(195)) or (inputs(247));
    layer0_outputs(8406) <= (inputs(17)) or (inputs(121));
    layer0_outputs(8407) <= inputs(175);
    layer0_outputs(8408) <= not((inputs(244)) or (inputs(181)));
    layer0_outputs(8409) <= '1';
    layer0_outputs(8410) <= (inputs(150)) and not (inputs(143));
    layer0_outputs(8411) <= not(inputs(41)) or (inputs(6));
    layer0_outputs(8412) <= not((inputs(18)) or (inputs(123)));
    layer0_outputs(8413) <= not(inputs(19));
    layer0_outputs(8414) <= not(inputs(95));
    layer0_outputs(8415) <= not((inputs(81)) and (inputs(140)));
    layer0_outputs(8416) <= (inputs(228)) and not (inputs(61));
    layer0_outputs(8417) <= (inputs(222)) or (inputs(164));
    layer0_outputs(8418) <= not(inputs(198));
    layer0_outputs(8419) <= not((inputs(5)) xor (inputs(222)));
    layer0_outputs(8420) <= not(inputs(107));
    layer0_outputs(8421) <= (inputs(217)) xor (inputs(200));
    layer0_outputs(8422) <= not((inputs(61)) or (inputs(144)));
    layer0_outputs(8423) <= '0';
    layer0_outputs(8424) <= not((inputs(32)) or (inputs(222)));
    layer0_outputs(8425) <= not((inputs(4)) or (inputs(155)));
    layer0_outputs(8426) <= not(inputs(117));
    layer0_outputs(8427) <= not((inputs(65)) and (inputs(187)));
    layer0_outputs(8428) <= not(inputs(160));
    layer0_outputs(8429) <= not(inputs(46)) or (inputs(0));
    layer0_outputs(8430) <= inputs(178);
    layer0_outputs(8431) <= not((inputs(0)) or (inputs(2)));
    layer0_outputs(8432) <= '1';
    layer0_outputs(8433) <= not(inputs(46));
    layer0_outputs(8434) <= (inputs(139)) or (inputs(100));
    layer0_outputs(8435) <= (inputs(14)) or (inputs(207));
    layer0_outputs(8436) <= not(inputs(161));
    layer0_outputs(8437) <= not((inputs(123)) xor (inputs(101)));
    layer0_outputs(8438) <= inputs(121);
    layer0_outputs(8439) <= inputs(2);
    layer0_outputs(8440) <= not(inputs(155)) or (inputs(241));
    layer0_outputs(8441) <= (inputs(172)) and not (inputs(207));
    layer0_outputs(8442) <= inputs(52);
    layer0_outputs(8443) <= (inputs(169)) and (inputs(185));
    layer0_outputs(8444) <= not(inputs(175)) or (inputs(186));
    layer0_outputs(8445) <= inputs(42);
    layer0_outputs(8446) <= (inputs(173)) or (inputs(175));
    layer0_outputs(8447) <= not(inputs(9));
    layer0_outputs(8448) <= (inputs(95)) xor (inputs(247));
    layer0_outputs(8449) <= not(inputs(60));
    layer0_outputs(8450) <= not(inputs(182));
    layer0_outputs(8451) <= not(inputs(85)) or (inputs(109));
    layer0_outputs(8452) <= not((inputs(4)) or (inputs(216)));
    layer0_outputs(8453) <= not(inputs(100));
    layer0_outputs(8454) <= not(inputs(117));
    layer0_outputs(8455) <= inputs(51);
    layer0_outputs(8456) <= not((inputs(48)) or (inputs(180)));
    layer0_outputs(8457) <= inputs(73);
    layer0_outputs(8458) <= (inputs(248)) and not (inputs(103));
    layer0_outputs(8459) <= not(inputs(123)) or (inputs(229));
    layer0_outputs(8460) <= '1';
    layer0_outputs(8461) <= (inputs(36)) and not (inputs(94));
    layer0_outputs(8462) <= not((inputs(31)) or (inputs(134)));
    layer0_outputs(8463) <= (inputs(112)) or (inputs(69));
    layer0_outputs(8464) <= not(inputs(95)) or (inputs(148));
    layer0_outputs(8465) <= not(inputs(178));
    layer0_outputs(8466) <= inputs(233);
    layer0_outputs(8467) <= not(inputs(151)) or (inputs(32));
    layer0_outputs(8468) <= (inputs(166)) and not (inputs(209));
    layer0_outputs(8469) <= (inputs(190)) or (inputs(9));
    layer0_outputs(8470) <= '1';
    layer0_outputs(8471) <= inputs(7);
    layer0_outputs(8472) <= not((inputs(226)) or (inputs(129)));
    layer0_outputs(8473) <= inputs(55);
    layer0_outputs(8474) <= not(inputs(166));
    layer0_outputs(8475) <= not(inputs(94));
    layer0_outputs(8476) <= not((inputs(150)) xor (inputs(3)));
    layer0_outputs(8477) <= (inputs(75)) xor (inputs(40));
    layer0_outputs(8478) <= not(inputs(41));
    layer0_outputs(8479) <= inputs(60);
    layer0_outputs(8480) <= inputs(253);
    layer0_outputs(8481) <= (inputs(100)) and not (inputs(231));
    layer0_outputs(8482) <= not(inputs(67)) or (inputs(166));
    layer0_outputs(8483) <= not((inputs(229)) xor (inputs(194)));
    layer0_outputs(8484) <= not(inputs(211));
    layer0_outputs(8485) <= (inputs(184)) and (inputs(249));
    layer0_outputs(8486) <= not(inputs(89));
    layer0_outputs(8487) <= (inputs(209)) or (inputs(71));
    layer0_outputs(8488) <= not(inputs(14)) or (inputs(76));
    layer0_outputs(8489) <= (inputs(161)) or (inputs(102));
    layer0_outputs(8490) <= '1';
    layer0_outputs(8491) <= (inputs(196)) and not (inputs(207));
    layer0_outputs(8492) <= not(inputs(113));
    layer0_outputs(8493) <= not(inputs(138));
    layer0_outputs(8494) <= not((inputs(152)) or (inputs(164)));
    layer0_outputs(8495) <= inputs(176);
    layer0_outputs(8496) <= inputs(5);
    layer0_outputs(8497) <= not(inputs(38)) or (inputs(178));
    layer0_outputs(8498) <= not(inputs(98)) or (inputs(12));
    layer0_outputs(8499) <= inputs(209);
    layer0_outputs(8500) <= inputs(115);
    layer0_outputs(8501) <= (inputs(143)) xor (inputs(246));
    layer0_outputs(8502) <= (inputs(196)) and not (inputs(15));
    layer0_outputs(8503) <= not(inputs(177));
    layer0_outputs(8504) <= inputs(202);
    layer0_outputs(8505) <= (inputs(219)) xor (inputs(225));
    layer0_outputs(8506) <= not((inputs(187)) or (inputs(88)));
    layer0_outputs(8507) <= not(inputs(134));
    layer0_outputs(8508) <= not(inputs(206)) or (inputs(79));
    layer0_outputs(8509) <= (inputs(108)) or (inputs(120));
    layer0_outputs(8510) <= not((inputs(85)) xor (inputs(131)));
    layer0_outputs(8511) <= (inputs(242)) or (inputs(176));
    layer0_outputs(8512) <= (inputs(235)) and not (inputs(80));
    layer0_outputs(8513) <= not((inputs(113)) or (inputs(43)));
    layer0_outputs(8514) <= not(inputs(211));
    layer0_outputs(8515) <= (inputs(12)) xor (inputs(56));
    layer0_outputs(8516) <= inputs(93);
    layer0_outputs(8517) <= not(inputs(20));
    layer0_outputs(8518) <= '1';
    layer0_outputs(8519) <= inputs(197);
    layer0_outputs(8520) <= not((inputs(59)) or (inputs(15)));
    layer0_outputs(8521) <= not((inputs(214)) or (inputs(230)));
    layer0_outputs(8522) <= '0';
    layer0_outputs(8523) <= not(inputs(39));
    layer0_outputs(8524) <= not(inputs(44));
    layer0_outputs(8525) <= inputs(24);
    layer0_outputs(8526) <= inputs(116);
    layer0_outputs(8527) <= not(inputs(23));
    layer0_outputs(8528) <= not(inputs(253));
    layer0_outputs(8529) <= not(inputs(128)) or (inputs(22));
    layer0_outputs(8530) <= not(inputs(113));
    layer0_outputs(8531) <= not(inputs(250));
    layer0_outputs(8532) <= not((inputs(75)) or (inputs(19)));
    layer0_outputs(8533) <= not((inputs(208)) or (inputs(210)));
    layer0_outputs(8534) <= inputs(252);
    layer0_outputs(8535) <= (inputs(71)) and not (inputs(122));
    layer0_outputs(8536) <= inputs(253);
    layer0_outputs(8537) <= (inputs(235)) xor (inputs(151));
    layer0_outputs(8538) <= not(inputs(162));
    layer0_outputs(8539) <= not((inputs(196)) xor (inputs(149)));
    layer0_outputs(8540) <= (inputs(195)) or (inputs(204));
    layer0_outputs(8541) <= (inputs(180)) and (inputs(244));
    layer0_outputs(8542) <= (inputs(177)) or (inputs(115));
    layer0_outputs(8543) <= (inputs(144)) xor (inputs(179));
    layer0_outputs(8544) <= inputs(14);
    layer0_outputs(8545) <= not((inputs(105)) and (inputs(84)));
    layer0_outputs(8546) <= (inputs(166)) and (inputs(221));
    layer0_outputs(8547) <= not(inputs(206));
    layer0_outputs(8548) <= (inputs(212)) and not (inputs(249));
    layer0_outputs(8549) <= inputs(79);
    layer0_outputs(8550) <= not(inputs(31));
    layer0_outputs(8551) <= (inputs(203)) or (inputs(67));
    layer0_outputs(8552) <= (inputs(46)) xor (inputs(61));
    layer0_outputs(8553) <= not((inputs(174)) or (inputs(34)));
    layer0_outputs(8554) <= not(inputs(228)) or (inputs(181));
    layer0_outputs(8555) <= '1';
    layer0_outputs(8556) <= (inputs(109)) or (inputs(84));
    layer0_outputs(8557) <= (inputs(181)) and not (inputs(50));
    layer0_outputs(8558) <= not(inputs(149));
    layer0_outputs(8559) <= (inputs(144)) or (inputs(12));
    layer0_outputs(8560) <= inputs(215);
    layer0_outputs(8561) <= not((inputs(248)) and (inputs(21)));
    layer0_outputs(8562) <= not(inputs(10));
    layer0_outputs(8563) <= not((inputs(45)) xor (inputs(131)));
    layer0_outputs(8564) <= not(inputs(219));
    layer0_outputs(8565) <= not(inputs(205)) or (inputs(99));
    layer0_outputs(8566) <= not(inputs(246));
    layer0_outputs(8567) <= (inputs(67)) or (inputs(75));
    layer0_outputs(8568) <= (inputs(120)) or (inputs(1));
    layer0_outputs(8569) <= not((inputs(71)) xor (inputs(8)));
    layer0_outputs(8570) <= (inputs(12)) or (inputs(36));
    layer0_outputs(8571) <= not((inputs(52)) or (inputs(64)));
    layer0_outputs(8572) <= not((inputs(120)) and (inputs(119)));
    layer0_outputs(8573) <= (inputs(56)) and (inputs(211));
    layer0_outputs(8574) <= inputs(151);
    layer0_outputs(8575) <= not((inputs(9)) or (inputs(195)));
    layer0_outputs(8576) <= not(inputs(116)) or (inputs(4));
    layer0_outputs(8577) <= not(inputs(122)) or (inputs(195));
    layer0_outputs(8578) <= inputs(196);
    layer0_outputs(8579) <= inputs(63);
    layer0_outputs(8580) <= inputs(203);
    layer0_outputs(8581) <= (inputs(85)) and (inputs(3));
    layer0_outputs(8582) <= not((inputs(53)) or (inputs(48)));
    layer0_outputs(8583) <= '1';
    layer0_outputs(8584) <= not(inputs(229));
    layer0_outputs(8585) <= not(inputs(137));
    layer0_outputs(8586) <= not(inputs(234));
    layer0_outputs(8587) <= not(inputs(12)) or (inputs(48));
    layer0_outputs(8588) <= not(inputs(122));
    layer0_outputs(8589) <= not((inputs(162)) or (inputs(107)));
    layer0_outputs(8590) <= not((inputs(121)) xor (inputs(17)));
    layer0_outputs(8591) <= not(inputs(225));
    layer0_outputs(8592) <= (inputs(57)) or (inputs(42));
    layer0_outputs(8593) <= (inputs(44)) xor (inputs(40));
    layer0_outputs(8594) <= not((inputs(227)) or (inputs(34)));
    layer0_outputs(8595) <= not(inputs(61)) or (inputs(206));
    layer0_outputs(8596) <= inputs(164);
    layer0_outputs(8597) <= not(inputs(247)) or (inputs(71));
    layer0_outputs(8598) <= (inputs(56)) and not (inputs(188));
    layer0_outputs(8599) <= not(inputs(149));
    layer0_outputs(8600) <= not((inputs(97)) xor (inputs(115)));
    layer0_outputs(8601) <= not(inputs(79));
    layer0_outputs(8602) <= (inputs(192)) xor (inputs(175));
    layer0_outputs(8603) <= not((inputs(107)) or (inputs(38)));
    layer0_outputs(8604) <= (inputs(162)) or (inputs(171));
    layer0_outputs(8605) <= inputs(99);
    layer0_outputs(8606) <= not((inputs(51)) xor (inputs(209)));
    layer0_outputs(8607) <= not(inputs(100)) or (inputs(227));
    layer0_outputs(8608) <= inputs(10);
    layer0_outputs(8609) <= not((inputs(108)) or (inputs(24)));
    layer0_outputs(8610) <= not(inputs(162)) or (inputs(76));
    layer0_outputs(8611) <= not((inputs(169)) or (inputs(164)));
    layer0_outputs(8612) <= '0';
    layer0_outputs(8613) <= inputs(102);
    layer0_outputs(8614) <= not(inputs(160)) or (inputs(241));
    layer0_outputs(8615) <= not(inputs(47)) or (inputs(28));
    layer0_outputs(8616) <= (inputs(19)) and not (inputs(35));
    layer0_outputs(8617) <= not(inputs(4));
    layer0_outputs(8618) <= not((inputs(67)) or (inputs(160)));
    layer0_outputs(8619) <= (inputs(210)) or (inputs(29));
    layer0_outputs(8620) <= (inputs(142)) or (inputs(186));
    layer0_outputs(8621) <= not(inputs(120));
    layer0_outputs(8622) <= not(inputs(183));
    layer0_outputs(8623) <= (inputs(125)) and not (inputs(140));
    layer0_outputs(8624) <= not((inputs(234)) xor (inputs(139)));
    layer0_outputs(8625) <= not(inputs(102));
    layer0_outputs(8626) <= not(inputs(220));
    layer0_outputs(8627) <= inputs(73);
    layer0_outputs(8628) <= inputs(58);
    layer0_outputs(8629) <= '0';
    layer0_outputs(8630) <= not((inputs(130)) or (inputs(159)));
    layer0_outputs(8631) <= not(inputs(227));
    layer0_outputs(8632) <= (inputs(78)) and not (inputs(199));
    layer0_outputs(8633) <= (inputs(184)) or (inputs(224));
    layer0_outputs(8634) <= (inputs(85)) or (inputs(149));
    layer0_outputs(8635) <= not(inputs(171)) or (inputs(158));
    layer0_outputs(8636) <= inputs(173);
    layer0_outputs(8637) <= not((inputs(190)) or (inputs(14)));
    layer0_outputs(8638) <= (inputs(180)) or (inputs(49));
    layer0_outputs(8639) <= '1';
    layer0_outputs(8640) <= (inputs(121)) and not (inputs(114));
    layer0_outputs(8641) <= not((inputs(204)) and (inputs(254)));
    layer0_outputs(8642) <= not(inputs(196)) or (inputs(92));
    layer0_outputs(8643) <= (inputs(240)) or (inputs(63));
    layer0_outputs(8644) <= inputs(133);
    layer0_outputs(8645) <= not((inputs(183)) and (inputs(111)));
    layer0_outputs(8646) <= not(inputs(99));
    layer0_outputs(8647) <= not((inputs(9)) xor (inputs(190)));
    layer0_outputs(8648) <= '0';
    layer0_outputs(8649) <= not((inputs(108)) or (inputs(175)));
    layer0_outputs(8650) <= not((inputs(84)) or (inputs(121)));
    layer0_outputs(8651) <= not(inputs(79)) or (inputs(8));
    layer0_outputs(8652) <= '1';
    layer0_outputs(8653) <= (inputs(2)) or (inputs(231));
    layer0_outputs(8654) <= (inputs(187)) and (inputs(226));
    layer0_outputs(8655) <= not((inputs(12)) and (inputs(230)));
    layer0_outputs(8656) <= inputs(148);
    layer0_outputs(8657) <= (inputs(21)) or (inputs(56));
    layer0_outputs(8658) <= not(inputs(179));
    layer0_outputs(8659) <= (inputs(232)) or (inputs(209));
    layer0_outputs(8660) <= not(inputs(174));
    layer0_outputs(8661) <= not((inputs(112)) or (inputs(225)));
    layer0_outputs(8662) <= not(inputs(100));
    layer0_outputs(8663) <= not(inputs(218));
    layer0_outputs(8664) <= (inputs(203)) and not (inputs(83));
    layer0_outputs(8665) <= inputs(56);
    layer0_outputs(8666) <= not(inputs(68));
    layer0_outputs(8667) <= (inputs(90)) and not (inputs(218));
    layer0_outputs(8668) <= (inputs(198)) or (inputs(115));
    layer0_outputs(8669) <= (inputs(60)) and not (inputs(12));
    layer0_outputs(8670) <= not((inputs(60)) or (inputs(184)));
    layer0_outputs(8671) <= not(inputs(214));
    layer0_outputs(8672) <= not((inputs(135)) or (inputs(208)));
    layer0_outputs(8673) <= not((inputs(22)) and (inputs(152)));
    layer0_outputs(8674) <= not(inputs(180));
    layer0_outputs(8675) <= '0';
    layer0_outputs(8676) <= not(inputs(218)) or (inputs(12));
    layer0_outputs(8677) <= (inputs(193)) or (inputs(192));
    layer0_outputs(8678) <= (inputs(253)) or (inputs(179));
    layer0_outputs(8679) <= (inputs(6)) and not (inputs(208));
    layer0_outputs(8680) <= (inputs(197)) or (inputs(49));
    layer0_outputs(8681) <= inputs(161);
    layer0_outputs(8682) <= not(inputs(125)) or (inputs(62));
    layer0_outputs(8683) <= (inputs(138)) or (inputs(145));
    layer0_outputs(8684) <= not(inputs(157));
    layer0_outputs(8685) <= inputs(171);
    layer0_outputs(8686) <= inputs(227);
    layer0_outputs(8687) <= not(inputs(9));
    layer0_outputs(8688) <= inputs(53);
    layer0_outputs(8689) <= not(inputs(97));
    layer0_outputs(8690) <= inputs(175);
    layer0_outputs(8691) <= inputs(134);
    layer0_outputs(8692) <= not((inputs(166)) or (inputs(113)));
    layer0_outputs(8693) <= not(inputs(198));
    layer0_outputs(8694) <= inputs(120);
    layer0_outputs(8695) <= '0';
    layer0_outputs(8696) <= not(inputs(200));
    layer0_outputs(8697) <= not(inputs(254));
    layer0_outputs(8698) <= (inputs(250)) or (inputs(116));
    layer0_outputs(8699) <= not(inputs(122));
    layer0_outputs(8700) <= not(inputs(240)) or (inputs(185));
    layer0_outputs(8701) <= (inputs(95)) or (inputs(148));
    layer0_outputs(8702) <= '1';
    layer0_outputs(8703) <= not((inputs(209)) and (inputs(239)));
    layer0_outputs(8704) <= not((inputs(202)) and (inputs(104)));
    layer0_outputs(8705) <= (inputs(5)) and not (inputs(224));
    layer0_outputs(8706) <= (inputs(172)) and not (inputs(14));
    layer0_outputs(8707) <= '1';
    layer0_outputs(8708) <= (inputs(155)) and not (inputs(239));
    layer0_outputs(8709) <= (inputs(110)) or (inputs(164));
    layer0_outputs(8710) <= not(inputs(139));
    layer0_outputs(8711) <= not((inputs(249)) xor (inputs(171)));
    layer0_outputs(8712) <= not(inputs(44)) or (inputs(122));
    layer0_outputs(8713) <= not(inputs(192));
    layer0_outputs(8714) <= (inputs(82)) or (inputs(164));
    layer0_outputs(8715) <= not(inputs(213));
    layer0_outputs(8716) <= not((inputs(242)) or (inputs(189)));
    layer0_outputs(8717) <= (inputs(170)) and not (inputs(112));
    layer0_outputs(8718) <= (inputs(127)) and not (inputs(216));
    layer0_outputs(8719) <= (inputs(106)) or (inputs(103));
    layer0_outputs(8720) <= (inputs(204)) or (inputs(179));
    layer0_outputs(8721) <= (inputs(89)) xor (inputs(136));
    layer0_outputs(8722) <= not(inputs(18)) or (inputs(111));
    layer0_outputs(8723) <= (inputs(1)) or (inputs(137));
    layer0_outputs(8724) <= not((inputs(58)) xor (inputs(37)));
    layer0_outputs(8725) <= (inputs(29)) or (inputs(177));
    layer0_outputs(8726) <= (inputs(229)) or (inputs(208));
    layer0_outputs(8727) <= (inputs(243)) xor (inputs(197));
    layer0_outputs(8728) <= (inputs(117)) xor (inputs(158));
    layer0_outputs(8729) <= (inputs(167)) and not (inputs(27));
    layer0_outputs(8730) <= not(inputs(105)) or (inputs(54));
    layer0_outputs(8731) <= inputs(26);
    layer0_outputs(8732) <= not((inputs(37)) or (inputs(39)));
    layer0_outputs(8733) <= (inputs(100)) and not (inputs(223));
    layer0_outputs(8734) <= not((inputs(98)) xor (inputs(50)));
    layer0_outputs(8735) <= not(inputs(193)) or (inputs(218));
    layer0_outputs(8736) <= not(inputs(186));
    layer0_outputs(8737) <= '0';
    layer0_outputs(8738) <= (inputs(239)) or (inputs(168));
    layer0_outputs(8739) <= (inputs(134)) and not (inputs(241));
    layer0_outputs(8740) <= not((inputs(209)) xor (inputs(205)));
    layer0_outputs(8741) <= (inputs(22)) or (inputs(160));
    layer0_outputs(8742) <= '1';
    layer0_outputs(8743) <= not(inputs(31)) or (inputs(241));
    layer0_outputs(8744) <= inputs(22);
    layer0_outputs(8745) <= not((inputs(7)) xor (inputs(16)));
    layer0_outputs(8746) <= not((inputs(195)) xor (inputs(103)));
    layer0_outputs(8747) <= not((inputs(218)) xor (inputs(250)));
    layer0_outputs(8748) <= inputs(254);
    layer0_outputs(8749) <= (inputs(84)) and not (inputs(190));
    layer0_outputs(8750) <= not((inputs(3)) or (inputs(24)));
    layer0_outputs(8751) <= (inputs(77)) and not (inputs(6));
    layer0_outputs(8752) <= not((inputs(249)) or (inputs(73)));
    layer0_outputs(8753) <= inputs(165);
    layer0_outputs(8754) <= (inputs(140)) and not (inputs(170));
    layer0_outputs(8755) <= not(inputs(139)) or (inputs(248));
    layer0_outputs(8756) <= (inputs(148)) and (inputs(9));
    layer0_outputs(8757) <= (inputs(157)) and not (inputs(49));
    layer0_outputs(8758) <= (inputs(129)) or (inputs(170));
    layer0_outputs(8759) <= not(inputs(212)) or (inputs(168));
    layer0_outputs(8760) <= not(inputs(231));
    layer0_outputs(8761) <= not((inputs(142)) and (inputs(189)));
    layer0_outputs(8762) <= not(inputs(85)) or (inputs(236));
    layer0_outputs(8763) <= inputs(230);
    layer0_outputs(8764) <= inputs(202);
    layer0_outputs(8765) <= not(inputs(85));
    layer0_outputs(8766) <= not((inputs(174)) or (inputs(171)));
    layer0_outputs(8767) <= not((inputs(103)) or (inputs(207)));
    layer0_outputs(8768) <= (inputs(1)) and (inputs(203));
    layer0_outputs(8769) <= inputs(110);
    layer0_outputs(8770) <= not(inputs(168));
    layer0_outputs(8771) <= (inputs(200)) and not (inputs(88));
    layer0_outputs(8772) <= not(inputs(136)) or (inputs(98));
    layer0_outputs(8773) <= not((inputs(109)) and (inputs(179)));
    layer0_outputs(8774) <= (inputs(16)) xor (inputs(77));
    layer0_outputs(8775) <= (inputs(148)) and not (inputs(173));
    layer0_outputs(8776) <= not((inputs(17)) xor (inputs(9)));
    layer0_outputs(8777) <= not(inputs(89)) or (inputs(173));
    layer0_outputs(8778) <= not(inputs(124));
    layer0_outputs(8779) <= not(inputs(76)) or (inputs(252));
    layer0_outputs(8780) <= inputs(89);
    layer0_outputs(8781) <= '0';
    layer0_outputs(8782) <= inputs(166);
    layer0_outputs(8783) <= not(inputs(147));
    layer0_outputs(8784) <= not(inputs(152)) or (inputs(48));
    layer0_outputs(8785) <= (inputs(149)) and not (inputs(59));
    layer0_outputs(8786) <= not(inputs(134)) or (inputs(76));
    layer0_outputs(8787) <= not((inputs(116)) or (inputs(196)));
    layer0_outputs(8788) <= not(inputs(206)) or (inputs(14));
    layer0_outputs(8789) <= (inputs(189)) and not (inputs(119));
    layer0_outputs(8790) <= not((inputs(157)) or (inputs(238)));
    layer0_outputs(8791) <= inputs(81);
    layer0_outputs(8792) <= inputs(179);
    layer0_outputs(8793) <= inputs(0);
    layer0_outputs(8794) <= inputs(106);
    layer0_outputs(8795) <= (inputs(201)) or (inputs(215));
    layer0_outputs(8796) <= (inputs(152)) and (inputs(144));
    layer0_outputs(8797) <= (inputs(194)) xor (inputs(208));
    layer0_outputs(8798) <= not(inputs(222));
    layer0_outputs(8799) <= not((inputs(96)) xor (inputs(126)));
    layer0_outputs(8800) <= not(inputs(11));
    layer0_outputs(8801) <= inputs(255);
    layer0_outputs(8802) <= (inputs(38)) or (inputs(61));
    layer0_outputs(8803) <= not((inputs(121)) xor (inputs(179)));
    layer0_outputs(8804) <= (inputs(193)) xor (inputs(38));
    layer0_outputs(8805) <= not(inputs(130));
    layer0_outputs(8806) <= not((inputs(206)) or (inputs(185)));
    layer0_outputs(8807) <= not((inputs(74)) and (inputs(241)));
    layer0_outputs(8808) <= '0';
    layer0_outputs(8809) <= (inputs(242)) and not (inputs(84));
    layer0_outputs(8810) <= not(inputs(146));
    layer0_outputs(8811) <= not((inputs(180)) or (inputs(188)));
    layer0_outputs(8812) <= (inputs(250)) or (inputs(128));
    layer0_outputs(8813) <= '1';
    layer0_outputs(8814) <= (inputs(139)) and not (inputs(212));
    layer0_outputs(8815) <= not(inputs(216)) or (inputs(78));
    layer0_outputs(8816) <= not(inputs(201)) or (inputs(4));
    layer0_outputs(8817) <= not(inputs(105));
    layer0_outputs(8818) <= inputs(56);
    layer0_outputs(8819) <= not((inputs(1)) and (inputs(83)));
    layer0_outputs(8820) <= inputs(36);
    layer0_outputs(8821) <= not(inputs(57));
    layer0_outputs(8822) <= not(inputs(199)) or (inputs(114));
    layer0_outputs(8823) <= (inputs(44)) or (inputs(245));
    layer0_outputs(8824) <= (inputs(155)) and not (inputs(65));
    layer0_outputs(8825) <= inputs(56);
    layer0_outputs(8826) <= not((inputs(205)) xor (inputs(241)));
    layer0_outputs(8827) <= not(inputs(22)) or (inputs(225));
    layer0_outputs(8828) <= inputs(52);
    layer0_outputs(8829) <= not(inputs(155)) or (inputs(46));
    layer0_outputs(8830) <= inputs(212);
    layer0_outputs(8831) <= (inputs(138)) and not (inputs(248));
    layer0_outputs(8832) <= not((inputs(48)) or (inputs(199)));
    layer0_outputs(8833) <= not(inputs(60));
    layer0_outputs(8834) <= '1';
    layer0_outputs(8835) <= (inputs(166)) and not (inputs(251));
    layer0_outputs(8836) <= inputs(234);
    layer0_outputs(8837) <= not(inputs(229)) or (inputs(60));
    layer0_outputs(8838) <= not((inputs(45)) and (inputs(216)));
    layer0_outputs(8839) <= not(inputs(168));
    layer0_outputs(8840) <= (inputs(149)) and not (inputs(16));
    layer0_outputs(8841) <= not((inputs(217)) or (inputs(96)));
    layer0_outputs(8842) <= not(inputs(52));
    layer0_outputs(8843) <= (inputs(57)) and not (inputs(49));
    layer0_outputs(8844) <= inputs(217);
    layer0_outputs(8845) <= inputs(92);
    layer0_outputs(8846) <= not(inputs(149));
    layer0_outputs(8847) <= (inputs(215)) and not (inputs(63));
    layer0_outputs(8848) <= '0';
    layer0_outputs(8849) <= (inputs(93)) or (inputs(46));
    layer0_outputs(8850) <= not(inputs(245));
    layer0_outputs(8851) <= (inputs(90)) or (inputs(102));
    layer0_outputs(8852) <= not(inputs(235));
    layer0_outputs(8853) <= not(inputs(60));
    layer0_outputs(8854) <= inputs(170);
    layer0_outputs(8855) <= not((inputs(146)) or (inputs(174)));
    layer0_outputs(8856) <= not(inputs(109)) or (inputs(147));
    layer0_outputs(8857) <= not(inputs(253));
    layer0_outputs(8858) <= not((inputs(10)) and (inputs(118)));
    layer0_outputs(8859) <= inputs(60);
    layer0_outputs(8860) <= not(inputs(58));
    layer0_outputs(8861) <= not(inputs(74));
    layer0_outputs(8862) <= (inputs(223)) xor (inputs(166));
    layer0_outputs(8863) <= (inputs(200)) and (inputs(202));
    layer0_outputs(8864) <= not((inputs(79)) or (inputs(107)));
    layer0_outputs(8865) <= not((inputs(62)) or (inputs(39)));
    layer0_outputs(8866) <= not(inputs(63)) or (inputs(248));
    layer0_outputs(8867) <= not((inputs(192)) or (inputs(35)));
    layer0_outputs(8868) <= not(inputs(218));
    layer0_outputs(8869) <= not(inputs(243)) or (inputs(203));
    layer0_outputs(8870) <= (inputs(101)) or (inputs(83));
    layer0_outputs(8871) <= '0';
    layer0_outputs(8872) <= not((inputs(227)) or (inputs(204)));
    layer0_outputs(8873) <= inputs(130);
    layer0_outputs(8874) <= inputs(229);
    layer0_outputs(8875) <= (inputs(67)) or (inputs(62));
    layer0_outputs(8876) <= inputs(182);
    layer0_outputs(8877) <= (inputs(176)) or (inputs(141));
    layer0_outputs(8878) <= not((inputs(117)) xor (inputs(153)));
    layer0_outputs(8879) <= not(inputs(6));
    layer0_outputs(8880) <= (inputs(185)) and (inputs(243));
    layer0_outputs(8881) <= not((inputs(49)) or (inputs(110)));
    layer0_outputs(8882) <= (inputs(79)) xor (inputs(76));
    layer0_outputs(8883) <= (inputs(249)) and not (inputs(253));
    layer0_outputs(8884) <= not(inputs(74));
    layer0_outputs(8885) <= not((inputs(80)) xor (inputs(11)));
    layer0_outputs(8886) <= (inputs(206)) and not (inputs(18));
    layer0_outputs(8887) <= inputs(1);
    layer0_outputs(8888) <= (inputs(181)) xor (inputs(182));
    layer0_outputs(8889) <= inputs(101);
    layer0_outputs(8890) <= '0';
    layer0_outputs(8891) <= inputs(154);
    layer0_outputs(8892) <= (inputs(59)) and not (inputs(192));
    layer0_outputs(8893) <= not((inputs(75)) and (inputs(218)));
    layer0_outputs(8894) <= inputs(194);
    layer0_outputs(8895) <= inputs(88);
    layer0_outputs(8896) <= not(inputs(77));
    layer0_outputs(8897) <= not(inputs(58));
    layer0_outputs(8898) <= (inputs(179)) and not (inputs(237));
    layer0_outputs(8899) <= not(inputs(57));
    layer0_outputs(8900) <= (inputs(73)) or (inputs(107));
    layer0_outputs(8901) <= (inputs(168)) and not (inputs(211));
    layer0_outputs(8902) <= not(inputs(154)) or (inputs(251));
    layer0_outputs(8903) <= not((inputs(7)) and (inputs(89)));
    layer0_outputs(8904) <= not(inputs(68));
    layer0_outputs(8905) <= not(inputs(56)) or (inputs(198));
    layer0_outputs(8906) <= (inputs(162)) or (inputs(155));
    layer0_outputs(8907) <= (inputs(124)) or (inputs(106));
    layer0_outputs(8908) <= '0';
    layer0_outputs(8909) <= inputs(102);
    layer0_outputs(8910) <= inputs(134);
    layer0_outputs(8911) <= '1';
    layer0_outputs(8912) <= (inputs(98)) and not (inputs(244));
    layer0_outputs(8913) <= (inputs(5)) or (inputs(216));
    layer0_outputs(8914) <= not(inputs(242)) or (inputs(34));
    layer0_outputs(8915) <= not(inputs(83)) or (inputs(191));
    layer0_outputs(8916) <= not(inputs(7)) or (inputs(209));
    layer0_outputs(8917) <= '0';
    layer0_outputs(8918) <= inputs(75);
    layer0_outputs(8919) <= (inputs(179)) or (inputs(111));
    layer0_outputs(8920) <= inputs(110);
    layer0_outputs(8921) <= not(inputs(190));
    layer0_outputs(8922) <= not(inputs(169));
    layer0_outputs(8923) <= not(inputs(92));
    layer0_outputs(8924) <= not(inputs(38)) or (inputs(143));
    layer0_outputs(8925) <= not((inputs(67)) or (inputs(176)));
    layer0_outputs(8926) <= inputs(87);
    layer0_outputs(8927) <= not(inputs(22)) or (inputs(15));
    layer0_outputs(8928) <= (inputs(88)) or (inputs(59));
    layer0_outputs(8929) <= (inputs(104)) xor (inputs(66));
    layer0_outputs(8930) <= inputs(12);
    layer0_outputs(8931) <= not(inputs(191));
    layer0_outputs(8932) <= not(inputs(214));
    layer0_outputs(8933) <= not(inputs(208));
    layer0_outputs(8934) <= not(inputs(18));
    layer0_outputs(8935) <= (inputs(19)) or (inputs(178));
    layer0_outputs(8936) <= '0';
    layer0_outputs(8937) <= (inputs(51)) and not (inputs(144));
    layer0_outputs(8938) <= not((inputs(106)) or (inputs(52)));
    layer0_outputs(8939) <= not((inputs(153)) or (inputs(207)));
    layer0_outputs(8940) <= not(inputs(206)) or (inputs(8));
    layer0_outputs(8941) <= (inputs(158)) and not (inputs(94));
    layer0_outputs(8942) <= (inputs(111)) or (inputs(196));
    layer0_outputs(8943) <= inputs(127);
    layer0_outputs(8944) <= not(inputs(50));
    layer0_outputs(8945) <= inputs(188);
    layer0_outputs(8946) <= '0';
    layer0_outputs(8947) <= inputs(43);
    layer0_outputs(8948) <= not(inputs(3)) or (inputs(172));
    layer0_outputs(8949) <= not((inputs(238)) and (inputs(13)));
    layer0_outputs(8950) <= not(inputs(79));
    layer0_outputs(8951) <= not(inputs(58));
    layer0_outputs(8952) <= (inputs(135)) or (inputs(241));
    layer0_outputs(8953) <= not((inputs(218)) and (inputs(208)));
    layer0_outputs(8954) <= not((inputs(239)) and (inputs(0)));
    layer0_outputs(8955) <= not((inputs(12)) xor (inputs(26)));
    layer0_outputs(8956) <= (inputs(158)) or (inputs(129));
    layer0_outputs(8957) <= inputs(100);
    layer0_outputs(8958) <= not(inputs(183));
    layer0_outputs(8959) <= inputs(114);
    layer0_outputs(8960) <= not(inputs(226));
    layer0_outputs(8961) <= (inputs(124)) and not (inputs(72));
    layer0_outputs(8962) <= not((inputs(29)) or (inputs(1)));
    layer0_outputs(8963) <= not(inputs(18));
    layer0_outputs(8964) <= inputs(167);
    layer0_outputs(8965) <= (inputs(194)) or (inputs(113));
    layer0_outputs(8966) <= not(inputs(152)) or (inputs(245));
    layer0_outputs(8967) <= (inputs(157)) and not (inputs(168));
    layer0_outputs(8968) <= not(inputs(179));
    layer0_outputs(8969) <= (inputs(121)) and not (inputs(86));
    layer0_outputs(8970) <= (inputs(44)) and not (inputs(145));
    layer0_outputs(8971) <= not((inputs(206)) and (inputs(35)));
    layer0_outputs(8972) <= not((inputs(28)) and (inputs(245)));
    layer0_outputs(8973) <= inputs(135);
    layer0_outputs(8974) <= (inputs(115)) or (inputs(114));
    layer0_outputs(8975) <= not(inputs(154));
    layer0_outputs(8976) <= inputs(58);
    layer0_outputs(8977) <= (inputs(247)) and not (inputs(183));
    layer0_outputs(8978) <= inputs(232);
    layer0_outputs(8979) <= not((inputs(103)) or (inputs(226)));
    layer0_outputs(8980) <= not((inputs(133)) xor (inputs(102)));
    layer0_outputs(8981) <= (inputs(29)) or (inputs(19));
    layer0_outputs(8982) <= (inputs(210)) or (inputs(98));
    layer0_outputs(8983) <= not((inputs(45)) or (inputs(34)));
    layer0_outputs(8984) <= not(inputs(139));
    layer0_outputs(8985) <= (inputs(208)) and (inputs(241));
    layer0_outputs(8986) <= not(inputs(250)) or (inputs(128));
    layer0_outputs(8987) <= not(inputs(61));
    layer0_outputs(8988) <= not((inputs(111)) xor (inputs(8)));
    layer0_outputs(8989) <= inputs(67);
    layer0_outputs(8990) <= inputs(222);
    layer0_outputs(8991) <= not((inputs(217)) and (inputs(216)));
    layer0_outputs(8992) <= (inputs(114)) or (inputs(1));
    layer0_outputs(8993) <= not(inputs(104));
    layer0_outputs(8994) <= inputs(117);
    layer0_outputs(8995) <= inputs(129);
    layer0_outputs(8996) <= (inputs(165)) xor (inputs(104));
    layer0_outputs(8997) <= not(inputs(98));
    layer0_outputs(8998) <= not(inputs(87)) or (inputs(176));
    layer0_outputs(8999) <= (inputs(226)) and (inputs(39));
    layer0_outputs(9000) <= (inputs(196)) or (inputs(143));
    layer0_outputs(9001) <= not(inputs(23));
    layer0_outputs(9002) <= (inputs(120)) and not (inputs(174));
    layer0_outputs(9003) <= inputs(88);
    layer0_outputs(9004) <= not(inputs(71));
    layer0_outputs(9005) <= not(inputs(219));
    layer0_outputs(9006) <= (inputs(13)) and (inputs(115));
    layer0_outputs(9007) <= (inputs(235)) and (inputs(202));
    layer0_outputs(9008) <= '0';
    layer0_outputs(9009) <= (inputs(184)) and not (inputs(41));
    layer0_outputs(9010) <= inputs(198);
    layer0_outputs(9011) <= not(inputs(236)) or (inputs(107));
    layer0_outputs(9012) <= (inputs(35)) and (inputs(33));
    layer0_outputs(9013) <= not(inputs(83));
    layer0_outputs(9014) <= not((inputs(73)) or (inputs(190)));
    layer0_outputs(9015) <= (inputs(132)) and (inputs(152));
    layer0_outputs(9016) <= not(inputs(82));
    layer0_outputs(9017) <= inputs(203);
    layer0_outputs(9018) <= not(inputs(28)) or (inputs(253));
    layer0_outputs(9019) <= inputs(233);
    layer0_outputs(9020) <= not(inputs(99));
    layer0_outputs(9021) <= not(inputs(232));
    layer0_outputs(9022) <= (inputs(116)) or (inputs(121));
    layer0_outputs(9023) <= not((inputs(227)) or (inputs(115)));
    layer0_outputs(9024) <= inputs(103);
    layer0_outputs(9025) <= not(inputs(192));
    layer0_outputs(9026) <= '0';
    layer0_outputs(9027) <= (inputs(166)) or (inputs(137));
    layer0_outputs(9028) <= not((inputs(172)) or (inputs(217)));
    layer0_outputs(9029) <= not(inputs(228));
    layer0_outputs(9030) <= not((inputs(59)) xor (inputs(44)));
    layer0_outputs(9031) <= '1';
    layer0_outputs(9032) <= not(inputs(132)) or (inputs(32));
    layer0_outputs(9033) <= not(inputs(49));
    layer0_outputs(9034) <= '0';
    layer0_outputs(9035) <= (inputs(70)) and not (inputs(65));
    layer0_outputs(9036) <= (inputs(190)) or (inputs(155));
    layer0_outputs(9037) <= not(inputs(1)) or (inputs(250));
    layer0_outputs(9038) <= not(inputs(170)) or (inputs(214));
    layer0_outputs(9039) <= inputs(98);
    layer0_outputs(9040) <= inputs(216);
    layer0_outputs(9041) <= not((inputs(16)) and (inputs(12)));
    layer0_outputs(9042) <= not(inputs(2)) or (inputs(177));
    layer0_outputs(9043) <= not(inputs(41)) or (inputs(46));
    layer0_outputs(9044) <= inputs(176);
    layer0_outputs(9045) <= not((inputs(167)) or (inputs(207)));
    layer0_outputs(9046) <= not(inputs(142));
    layer0_outputs(9047) <= inputs(229);
    layer0_outputs(9048) <= (inputs(51)) or (inputs(80));
    layer0_outputs(9049) <= inputs(25);
    layer0_outputs(9050) <= not(inputs(189));
    layer0_outputs(9051) <= inputs(221);
    layer0_outputs(9052) <= (inputs(6)) or (inputs(18));
    layer0_outputs(9053) <= (inputs(145)) or (inputs(143));
    layer0_outputs(9054) <= not(inputs(197)) or (inputs(238));
    layer0_outputs(9055) <= not((inputs(34)) or (inputs(182)));
    layer0_outputs(9056) <= not(inputs(214));
    layer0_outputs(9057) <= (inputs(100)) and not (inputs(49));
    layer0_outputs(9058) <= inputs(27);
    layer0_outputs(9059) <= (inputs(184)) xor (inputs(119));
    layer0_outputs(9060) <= (inputs(29)) xor (inputs(47));
    layer0_outputs(9061) <= not(inputs(6));
    layer0_outputs(9062) <= (inputs(153)) or (inputs(24));
    layer0_outputs(9063) <= inputs(15);
    layer0_outputs(9064) <= '1';
    layer0_outputs(9065) <= not(inputs(24)) or (inputs(217));
    layer0_outputs(9066) <= (inputs(167)) or (inputs(254));
    layer0_outputs(9067) <= inputs(124);
    layer0_outputs(9068) <= inputs(118);
    layer0_outputs(9069) <= not(inputs(198));
    layer0_outputs(9070) <= (inputs(26)) and not (inputs(195));
    layer0_outputs(9071) <= not((inputs(78)) or (inputs(252)));
    layer0_outputs(9072) <= (inputs(208)) or (inputs(174));
    layer0_outputs(9073) <= inputs(81);
    layer0_outputs(9074) <= not(inputs(179));
    layer0_outputs(9075) <= '1';
    layer0_outputs(9076) <= (inputs(187)) and (inputs(184));
    layer0_outputs(9077) <= (inputs(135)) and not (inputs(5));
    layer0_outputs(9078) <= not(inputs(112)) or (inputs(54));
    layer0_outputs(9079) <= not(inputs(63)) or (inputs(16));
    layer0_outputs(9080) <= not((inputs(136)) or (inputs(80)));
    layer0_outputs(9081) <= '0';
    layer0_outputs(9082) <= not(inputs(84));
    layer0_outputs(9083) <= not(inputs(51)) or (inputs(198));
    layer0_outputs(9084) <= not(inputs(195));
    layer0_outputs(9085) <= inputs(176);
    layer0_outputs(9086) <= inputs(108);
    layer0_outputs(9087) <= not(inputs(118));
    layer0_outputs(9088) <= inputs(166);
    layer0_outputs(9089) <= not(inputs(179)) or (inputs(167));
    layer0_outputs(9090) <= not((inputs(103)) or (inputs(226)));
    layer0_outputs(9091) <= (inputs(119)) and not (inputs(82));
    layer0_outputs(9092) <= not(inputs(205)) or (inputs(191));
    layer0_outputs(9093) <= inputs(179);
    layer0_outputs(9094) <= not((inputs(86)) or (inputs(255)));
    layer0_outputs(9095) <= (inputs(202)) and not (inputs(146));
    layer0_outputs(9096) <= inputs(81);
    layer0_outputs(9097) <= not(inputs(37)) or (inputs(229));
    layer0_outputs(9098) <= not((inputs(120)) xor (inputs(174)));
    layer0_outputs(9099) <= not(inputs(6));
    layer0_outputs(9100) <= (inputs(9)) and (inputs(202));
    layer0_outputs(9101) <= not(inputs(246)) or (inputs(35));
    layer0_outputs(9102) <= (inputs(151)) and not (inputs(67));
    layer0_outputs(9103) <= inputs(243);
    layer0_outputs(9104) <= (inputs(164)) and not (inputs(185));
    layer0_outputs(9105) <= not(inputs(157)) or (inputs(15));
    layer0_outputs(9106) <= not(inputs(165));
    layer0_outputs(9107) <= (inputs(79)) and not (inputs(29));
    layer0_outputs(9108) <= not(inputs(119)) or (inputs(186));
    layer0_outputs(9109) <= (inputs(62)) and (inputs(195));
    layer0_outputs(9110) <= not((inputs(37)) or (inputs(56)));
    layer0_outputs(9111) <= inputs(21);
    layer0_outputs(9112) <= not(inputs(93)) or (inputs(203));
    layer0_outputs(9113) <= inputs(163);
    layer0_outputs(9114) <= not(inputs(118));
    layer0_outputs(9115) <= not((inputs(103)) or (inputs(5)));
    layer0_outputs(9116) <= inputs(107);
    layer0_outputs(9117) <= (inputs(157)) and (inputs(20));
    layer0_outputs(9118) <= inputs(167);
    layer0_outputs(9119) <= (inputs(163)) or (inputs(159));
    layer0_outputs(9120) <= not(inputs(155));
    layer0_outputs(9121) <= inputs(85);
    layer0_outputs(9122) <= (inputs(4)) and not (inputs(251));
    layer0_outputs(9123) <= (inputs(214)) xor (inputs(213));
    layer0_outputs(9124) <= not(inputs(169)) or (inputs(39));
    layer0_outputs(9125) <= inputs(26);
    layer0_outputs(9126) <= '0';
    layer0_outputs(9127) <= (inputs(54)) and not (inputs(96));
    layer0_outputs(9128) <= not(inputs(246));
    layer0_outputs(9129) <= (inputs(76)) and not (inputs(161));
    layer0_outputs(9130) <= (inputs(20)) and not (inputs(145));
    layer0_outputs(9131) <= inputs(124);
    layer0_outputs(9132) <= inputs(233);
    layer0_outputs(9133) <= (inputs(132)) and (inputs(92));
    layer0_outputs(9134) <= (inputs(152)) and not (inputs(204));
    layer0_outputs(9135) <= inputs(129);
    layer0_outputs(9136) <= inputs(98);
    layer0_outputs(9137) <= (inputs(181)) and (inputs(9));
    layer0_outputs(9138) <= (inputs(83)) and (inputs(43));
    layer0_outputs(9139) <= (inputs(71)) and not (inputs(222));
    layer0_outputs(9140) <= not((inputs(46)) and (inputs(77)));
    layer0_outputs(9141) <= not(inputs(101)) or (inputs(77));
    layer0_outputs(9142) <= (inputs(164)) xor (inputs(239));
    layer0_outputs(9143) <= not(inputs(158));
    layer0_outputs(9144) <= inputs(150);
    layer0_outputs(9145) <= not(inputs(85));
    layer0_outputs(9146) <= not(inputs(85));
    layer0_outputs(9147) <= inputs(61);
    layer0_outputs(9148) <= not(inputs(23)) or (inputs(188));
    layer0_outputs(9149) <= (inputs(155)) and (inputs(73));
    layer0_outputs(9150) <= (inputs(71)) and not (inputs(64));
    layer0_outputs(9151) <= not(inputs(147)) or (inputs(237));
    layer0_outputs(9152) <= inputs(97);
    layer0_outputs(9153) <= not((inputs(180)) or (inputs(164)));
    layer0_outputs(9154) <= not((inputs(64)) xor (inputs(26)));
    layer0_outputs(9155) <= (inputs(44)) and (inputs(75));
    layer0_outputs(9156) <= (inputs(181)) xor (inputs(211));
    layer0_outputs(9157) <= (inputs(36)) and (inputs(27));
    layer0_outputs(9158) <= inputs(105);
    layer0_outputs(9159) <= not(inputs(4)) or (inputs(179));
    layer0_outputs(9160) <= not((inputs(6)) xor (inputs(195)));
    layer0_outputs(9161) <= not(inputs(99)) or (inputs(0));
    layer0_outputs(9162) <= (inputs(229)) and not (inputs(66));
    layer0_outputs(9163) <= (inputs(160)) or (inputs(84));
    layer0_outputs(9164) <= not((inputs(134)) xor (inputs(225)));
    layer0_outputs(9165) <= not(inputs(107)) or (inputs(211));
    layer0_outputs(9166) <= not((inputs(198)) or (inputs(80)));
    layer0_outputs(9167) <= not(inputs(161));
    layer0_outputs(9168) <= not((inputs(125)) or (inputs(205)));
    layer0_outputs(9169) <= not(inputs(93));
    layer0_outputs(9170) <= (inputs(129)) xor (inputs(164));
    layer0_outputs(9171) <= not((inputs(104)) or (inputs(214)));
    layer0_outputs(9172) <= (inputs(184)) and (inputs(253));
    layer0_outputs(9173) <= not((inputs(63)) xor (inputs(157)));
    layer0_outputs(9174) <= not(inputs(219)) or (inputs(249));
    layer0_outputs(9175) <= (inputs(3)) and not (inputs(47));
    layer0_outputs(9176) <= not((inputs(171)) and (inputs(42)));
    layer0_outputs(9177) <= not(inputs(221));
    layer0_outputs(9178) <= not(inputs(242)) or (inputs(97));
    layer0_outputs(9179) <= (inputs(189)) and not (inputs(178));
    layer0_outputs(9180) <= not(inputs(128)) or (inputs(251));
    layer0_outputs(9181) <= (inputs(58)) and (inputs(192));
    layer0_outputs(9182) <= (inputs(232)) xor (inputs(217));
    layer0_outputs(9183) <= inputs(82);
    layer0_outputs(9184) <= not((inputs(106)) or (inputs(255)));
    layer0_outputs(9185) <= not((inputs(169)) or (inputs(236)));
    layer0_outputs(9186) <= inputs(218);
    layer0_outputs(9187) <= '0';
    layer0_outputs(9188) <= not(inputs(196));
    layer0_outputs(9189) <= (inputs(11)) xor (inputs(76));
    layer0_outputs(9190) <= not(inputs(79));
    layer0_outputs(9191) <= not(inputs(141));
    layer0_outputs(9192) <= (inputs(93)) or (inputs(73));
    layer0_outputs(9193) <= not(inputs(167));
    layer0_outputs(9194) <= '0';
    layer0_outputs(9195) <= not((inputs(78)) or (inputs(44)));
    layer0_outputs(9196) <= not(inputs(210));
    layer0_outputs(9197) <= not((inputs(167)) xor (inputs(148)));
    layer0_outputs(9198) <= '0';
    layer0_outputs(9199) <= (inputs(99)) and not (inputs(56));
    layer0_outputs(9200) <= '1';
    layer0_outputs(9201) <= '1';
    layer0_outputs(9202) <= not((inputs(26)) or (inputs(58)));
    layer0_outputs(9203) <= inputs(199);
    layer0_outputs(9204) <= '1';
    layer0_outputs(9205) <= not(inputs(0)) or (inputs(242));
    layer0_outputs(9206) <= not((inputs(202)) or (inputs(129)));
    layer0_outputs(9207) <= (inputs(169)) and not (inputs(3));
    layer0_outputs(9208) <= (inputs(0)) and not (inputs(93));
    layer0_outputs(9209) <= (inputs(116)) and not (inputs(209));
    layer0_outputs(9210) <= not((inputs(186)) and (inputs(230)));
    layer0_outputs(9211) <= not(inputs(30)) or (inputs(42));
    layer0_outputs(9212) <= not((inputs(116)) or (inputs(142)));
    layer0_outputs(9213) <= (inputs(25)) and not (inputs(4));
    layer0_outputs(9214) <= not(inputs(177));
    layer0_outputs(9215) <= not(inputs(202));
    layer0_outputs(9216) <= not(inputs(166)) or (inputs(214));
    layer0_outputs(9217) <= not(inputs(22));
    layer0_outputs(9218) <= inputs(104);
    layer0_outputs(9219) <= (inputs(31)) and not (inputs(63));
    layer0_outputs(9220) <= (inputs(90)) xor (inputs(57));
    layer0_outputs(9221) <= not(inputs(41));
    layer0_outputs(9222) <= not(inputs(74)) or (inputs(49));
    layer0_outputs(9223) <= not((inputs(33)) or (inputs(110)));
    layer0_outputs(9224) <= inputs(115);
    layer0_outputs(9225) <= inputs(105);
    layer0_outputs(9226) <= not(inputs(230));
    layer0_outputs(9227) <= not(inputs(17));
    layer0_outputs(9228) <= not(inputs(20));
    layer0_outputs(9229) <= (inputs(81)) and not (inputs(106));
    layer0_outputs(9230) <= (inputs(138)) xor (inputs(218));
    layer0_outputs(9231) <= not(inputs(213)) or (inputs(98));
    layer0_outputs(9232) <= inputs(73);
    layer0_outputs(9233) <= inputs(177);
    layer0_outputs(9234) <= not(inputs(197));
    layer0_outputs(9235) <= inputs(233);
    layer0_outputs(9236) <= not(inputs(12)) or (inputs(197));
    layer0_outputs(9237) <= (inputs(190)) xor (inputs(143));
    layer0_outputs(9238) <= inputs(152);
    layer0_outputs(9239) <= not((inputs(54)) xor (inputs(22)));
    layer0_outputs(9240) <= not(inputs(172)) or (inputs(30));
    layer0_outputs(9241) <= (inputs(124)) xor (inputs(7));
    layer0_outputs(9242) <= not(inputs(55));
    layer0_outputs(9243) <= inputs(143);
    layer0_outputs(9244) <= (inputs(252)) or (inputs(114));
    layer0_outputs(9245) <= '0';
    layer0_outputs(9246) <= not(inputs(249));
    layer0_outputs(9247) <= (inputs(180)) and not (inputs(113));
    layer0_outputs(9248) <= not(inputs(125));
    layer0_outputs(9249) <= not(inputs(211));
    layer0_outputs(9250) <= (inputs(92)) or (inputs(90));
    layer0_outputs(9251) <= not(inputs(228));
    layer0_outputs(9252) <= not((inputs(162)) xor (inputs(118)));
    layer0_outputs(9253) <= not(inputs(131));
    layer0_outputs(9254) <= not(inputs(7)) or (inputs(53));
    layer0_outputs(9255) <= (inputs(84)) or (inputs(10));
    layer0_outputs(9256) <= not(inputs(249));
    layer0_outputs(9257) <= not((inputs(90)) xor (inputs(225)));
    layer0_outputs(9258) <= not((inputs(233)) or (inputs(236)));
    layer0_outputs(9259) <= not(inputs(44)) or (inputs(116));
    layer0_outputs(9260) <= '1';
    layer0_outputs(9261) <= not((inputs(54)) or (inputs(11)));
    layer0_outputs(9262) <= (inputs(141)) or (inputs(234));
    layer0_outputs(9263) <= not(inputs(37));
    layer0_outputs(9264) <= not(inputs(144));
    layer0_outputs(9265) <= '1';
    layer0_outputs(9266) <= (inputs(234)) and not (inputs(137));
    layer0_outputs(9267) <= not((inputs(124)) xor (inputs(95)));
    layer0_outputs(9268) <= not(inputs(124)) or (inputs(65));
    layer0_outputs(9269) <= inputs(32);
    layer0_outputs(9270) <= not(inputs(111));
    layer0_outputs(9271) <= (inputs(61)) xor (inputs(33));
    layer0_outputs(9272) <= (inputs(190)) xor (inputs(93));
    layer0_outputs(9273) <= (inputs(97)) and (inputs(146));
    layer0_outputs(9274) <= (inputs(195)) or (inputs(232));
    layer0_outputs(9275) <= not((inputs(63)) or (inputs(235)));
    layer0_outputs(9276) <= not(inputs(174));
    layer0_outputs(9277) <= not(inputs(189));
    layer0_outputs(9278) <= not(inputs(229)) or (inputs(20));
    layer0_outputs(9279) <= not((inputs(218)) or (inputs(161)));
    layer0_outputs(9280) <= inputs(54);
    layer0_outputs(9281) <= not((inputs(99)) xor (inputs(183)));
    layer0_outputs(9282) <= (inputs(183)) and not (inputs(60));
    layer0_outputs(9283) <= inputs(231);
    layer0_outputs(9284) <= not((inputs(26)) and (inputs(146)));
    layer0_outputs(9285) <= not(inputs(161));
    layer0_outputs(9286) <= (inputs(94)) and not (inputs(50));
    layer0_outputs(9287) <= inputs(95);
    layer0_outputs(9288) <= not(inputs(44));
    layer0_outputs(9289) <= (inputs(220)) or (inputs(231));
    layer0_outputs(9290) <= not(inputs(138));
    layer0_outputs(9291) <= (inputs(49)) and not (inputs(113));
    layer0_outputs(9292) <= (inputs(181)) or (inputs(8));
    layer0_outputs(9293) <= inputs(201);
    layer0_outputs(9294) <= (inputs(223)) xor (inputs(156));
    layer0_outputs(9295) <= not(inputs(232)) or (inputs(67));
    layer0_outputs(9296) <= not((inputs(182)) xor (inputs(216)));
    layer0_outputs(9297) <= not(inputs(166));
    layer0_outputs(9298) <= not(inputs(226)) or (inputs(108));
    layer0_outputs(9299) <= inputs(110);
    layer0_outputs(9300) <= inputs(248);
    layer0_outputs(9301) <= not(inputs(3));
    layer0_outputs(9302) <= '0';
    layer0_outputs(9303) <= (inputs(253)) and not (inputs(50));
    layer0_outputs(9304) <= not(inputs(23));
    layer0_outputs(9305) <= not(inputs(34)) or (inputs(252));
    layer0_outputs(9306) <= (inputs(64)) or (inputs(24));
    layer0_outputs(9307) <= (inputs(30)) or (inputs(159));
    layer0_outputs(9308) <= (inputs(79)) and not (inputs(66));
    layer0_outputs(9309) <= inputs(166);
    layer0_outputs(9310) <= not(inputs(73)) or (inputs(154));
    layer0_outputs(9311) <= not(inputs(138)) or (inputs(2));
    layer0_outputs(9312) <= (inputs(48)) and not (inputs(132));
    layer0_outputs(9313) <= not(inputs(227));
    layer0_outputs(9314) <= not((inputs(113)) or (inputs(9)));
    layer0_outputs(9315) <= not((inputs(137)) or (inputs(67)));
    layer0_outputs(9316) <= (inputs(79)) xor (inputs(179));
    layer0_outputs(9317) <= not((inputs(197)) or (inputs(231)));
    layer0_outputs(9318) <= (inputs(198)) and not (inputs(64));
    layer0_outputs(9319) <= not(inputs(210));
    layer0_outputs(9320) <= '0';
    layer0_outputs(9321) <= not((inputs(239)) xor (inputs(222)));
    layer0_outputs(9322) <= not(inputs(62)) or (inputs(33));
    layer0_outputs(9323) <= not((inputs(96)) xor (inputs(247)));
    layer0_outputs(9324) <= not(inputs(164)) or (inputs(156));
    layer0_outputs(9325) <= not(inputs(130));
    layer0_outputs(9326) <= (inputs(224)) or (inputs(63));
    layer0_outputs(9327) <= inputs(29);
    layer0_outputs(9328) <= (inputs(73)) and (inputs(166));
    layer0_outputs(9329) <= inputs(140);
    layer0_outputs(9330) <= not((inputs(132)) and (inputs(218)));
    layer0_outputs(9331) <= not(inputs(202));
    layer0_outputs(9332) <= not(inputs(241)) or (inputs(244));
    layer0_outputs(9333) <= not((inputs(11)) xor (inputs(42)));
    layer0_outputs(9334) <= not(inputs(123));
    layer0_outputs(9335) <= (inputs(64)) xor (inputs(23));
    layer0_outputs(9336) <= (inputs(104)) or (inputs(46));
    layer0_outputs(9337) <= not((inputs(235)) xor (inputs(229)));
    layer0_outputs(9338) <= not((inputs(151)) or (inputs(251)));
    layer0_outputs(9339) <= not((inputs(124)) or (inputs(139)));
    layer0_outputs(9340) <= not((inputs(203)) or (inputs(231)));
    layer0_outputs(9341) <= (inputs(18)) and not (inputs(107));
    layer0_outputs(9342) <= (inputs(167)) and not (inputs(13));
    layer0_outputs(9343) <= not((inputs(235)) xor (inputs(186)));
    layer0_outputs(9344) <= not((inputs(65)) and (inputs(245)));
    layer0_outputs(9345) <= (inputs(118)) and not (inputs(70));
    layer0_outputs(9346) <= (inputs(199)) and not (inputs(77));
    layer0_outputs(9347) <= not((inputs(24)) xor (inputs(91)));
    layer0_outputs(9348) <= inputs(3);
    layer0_outputs(9349) <= not((inputs(251)) or (inputs(112)));
    layer0_outputs(9350) <= (inputs(247)) or (inputs(243));
    layer0_outputs(9351) <= not((inputs(15)) or (inputs(121)));
    layer0_outputs(9352) <= (inputs(253)) or (inputs(135));
    layer0_outputs(9353) <= (inputs(19)) and not (inputs(223));
    layer0_outputs(9354) <= not((inputs(93)) xor (inputs(75)));
    layer0_outputs(9355) <= inputs(213);
    layer0_outputs(9356) <= inputs(74);
    layer0_outputs(9357) <= inputs(61);
    layer0_outputs(9358) <= not((inputs(175)) or (inputs(218)));
    layer0_outputs(9359) <= (inputs(147)) or (inputs(132));
    layer0_outputs(9360) <= inputs(145);
    layer0_outputs(9361) <= not((inputs(163)) and (inputs(18)));
    layer0_outputs(9362) <= not(inputs(121));
    layer0_outputs(9363) <= not((inputs(108)) or (inputs(106)));
    layer0_outputs(9364) <= '0';
    layer0_outputs(9365) <= not(inputs(8));
    layer0_outputs(9366) <= not(inputs(98));
    layer0_outputs(9367) <= (inputs(145)) or (inputs(217));
    layer0_outputs(9368) <= not((inputs(158)) xor (inputs(204)));
    layer0_outputs(9369) <= inputs(198);
    layer0_outputs(9370) <= not(inputs(201));
    layer0_outputs(9371) <= not(inputs(141)) or (inputs(248));
    layer0_outputs(9372) <= not(inputs(171)) or (inputs(14));
    layer0_outputs(9373) <= (inputs(192)) and not (inputs(98));
    layer0_outputs(9374) <= not(inputs(76));
    layer0_outputs(9375) <= (inputs(42)) and (inputs(79));
    layer0_outputs(9376) <= inputs(181);
    layer0_outputs(9377) <= not(inputs(232));
    layer0_outputs(9378) <= not((inputs(201)) or (inputs(225)));
    layer0_outputs(9379) <= inputs(94);
    layer0_outputs(9380) <= (inputs(61)) and not (inputs(113));
    layer0_outputs(9381) <= (inputs(207)) and not (inputs(16));
    layer0_outputs(9382) <= not((inputs(175)) or (inputs(144)));
    layer0_outputs(9383) <= not(inputs(106)) or (inputs(68));
    layer0_outputs(9384) <= '1';
    layer0_outputs(9385) <= (inputs(18)) and (inputs(30));
    layer0_outputs(9386) <= '0';
    layer0_outputs(9387) <= not(inputs(38)) or (inputs(148));
    layer0_outputs(9388) <= not(inputs(117));
    layer0_outputs(9389) <= not((inputs(217)) or (inputs(18)));
    layer0_outputs(9390) <= not((inputs(22)) xor (inputs(55)));
    layer0_outputs(9391) <= (inputs(134)) and not (inputs(225));
    layer0_outputs(9392) <= (inputs(148)) or (inputs(235));
    layer0_outputs(9393) <= not(inputs(249));
    layer0_outputs(9394) <= not(inputs(205)) or (inputs(78));
    layer0_outputs(9395) <= (inputs(107)) and not (inputs(158));
    layer0_outputs(9396) <= inputs(198);
    layer0_outputs(9397) <= not(inputs(206));
    layer0_outputs(9398) <= not(inputs(186)) or (inputs(113));
    layer0_outputs(9399) <= not(inputs(168));
    layer0_outputs(9400) <= not(inputs(94));
    layer0_outputs(9401) <= not(inputs(21));
    layer0_outputs(9402) <= not(inputs(245));
    layer0_outputs(9403) <= not((inputs(33)) or (inputs(23)));
    layer0_outputs(9404) <= '1';
    layer0_outputs(9405) <= not((inputs(165)) xor (inputs(130)));
    layer0_outputs(9406) <= (inputs(16)) and not (inputs(159));
    layer0_outputs(9407) <= not(inputs(125));
    layer0_outputs(9408) <= (inputs(33)) xor (inputs(142));
    layer0_outputs(9409) <= not((inputs(41)) or (inputs(83)));
    layer0_outputs(9410) <= inputs(130);
    layer0_outputs(9411) <= inputs(27);
    layer0_outputs(9412) <= (inputs(95)) and (inputs(123));
    layer0_outputs(9413) <= not((inputs(32)) or (inputs(224)));
    layer0_outputs(9414) <= (inputs(21)) and not (inputs(85));
    layer0_outputs(9415) <= '0';
    layer0_outputs(9416) <= not(inputs(6));
    layer0_outputs(9417) <= inputs(7);
    layer0_outputs(9418) <= (inputs(159)) or (inputs(248));
    layer0_outputs(9419) <= not(inputs(244)) or (inputs(8));
    layer0_outputs(9420) <= inputs(77);
    layer0_outputs(9421) <= not(inputs(94));
    layer0_outputs(9422) <= (inputs(15)) and not (inputs(7));
    layer0_outputs(9423) <= (inputs(164)) or (inputs(82));
    layer0_outputs(9424) <= not(inputs(20)) or (inputs(22));
    layer0_outputs(9425) <= not(inputs(55));
    layer0_outputs(9426) <= not(inputs(231));
    layer0_outputs(9427) <= not(inputs(163));
    layer0_outputs(9428) <= not(inputs(227)) or (inputs(16));
    layer0_outputs(9429) <= inputs(23);
    layer0_outputs(9430) <= not((inputs(91)) or (inputs(125)));
    layer0_outputs(9431) <= not(inputs(227));
    layer0_outputs(9432) <= not((inputs(234)) xor (inputs(42)));
    layer0_outputs(9433) <= (inputs(52)) xor (inputs(86));
    layer0_outputs(9434) <= (inputs(144)) and (inputs(115));
    layer0_outputs(9435) <= (inputs(18)) or (inputs(160));
    layer0_outputs(9436) <= inputs(25);
    layer0_outputs(9437) <= '0';
    layer0_outputs(9438) <= inputs(228);
    layer0_outputs(9439) <= (inputs(168)) and not (inputs(156));
    layer0_outputs(9440) <= not((inputs(98)) or (inputs(157)));
    layer0_outputs(9441) <= not(inputs(165));
    layer0_outputs(9442) <= (inputs(169)) or (inputs(33));
    layer0_outputs(9443) <= not(inputs(214));
    layer0_outputs(9444) <= (inputs(106)) and not (inputs(129));
    layer0_outputs(9445) <= not(inputs(114));
    layer0_outputs(9446) <= (inputs(150)) and not (inputs(196));
    layer0_outputs(9447) <= not(inputs(187));
    layer0_outputs(9448) <= not(inputs(59));
    layer0_outputs(9449) <= not(inputs(76));
    layer0_outputs(9450) <= (inputs(142)) and not (inputs(207));
    layer0_outputs(9451) <= (inputs(158)) or (inputs(33));
    layer0_outputs(9452) <= (inputs(149)) and not (inputs(255));
    layer0_outputs(9453) <= not(inputs(133));
    layer0_outputs(9454) <= inputs(58);
    layer0_outputs(9455) <= not((inputs(105)) or (inputs(135)));
    layer0_outputs(9456) <= not((inputs(238)) or (inputs(221)));
    layer0_outputs(9457) <= (inputs(125)) and not (inputs(254));
    layer0_outputs(9458) <= (inputs(175)) or (inputs(227));
    layer0_outputs(9459) <= inputs(66);
    layer0_outputs(9460) <= not(inputs(64));
    layer0_outputs(9461) <= not(inputs(148)) or (inputs(97));
    layer0_outputs(9462) <= (inputs(4)) or (inputs(131));
    layer0_outputs(9463) <= '1';
    layer0_outputs(9464) <= not(inputs(59));
    layer0_outputs(9465) <= not((inputs(254)) or (inputs(92)));
    layer0_outputs(9466) <= inputs(190);
    layer0_outputs(9467) <= inputs(166);
    layer0_outputs(9468) <= inputs(255);
    layer0_outputs(9469) <= not(inputs(188));
    layer0_outputs(9470) <= inputs(73);
    layer0_outputs(9471) <= not(inputs(229)) or (inputs(17));
    layer0_outputs(9472) <= not(inputs(230));
    layer0_outputs(9473) <= not(inputs(237));
    layer0_outputs(9474) <= not(inputs(157)) or (inputs(183));
    layer0_outputs(9475) <= not((inputs(68)) or (inputs(195)));
    layer0_outputs(9476) <= not((inputs(31)) or (inputs(124)));
    layer0_outputs(9477) <= (inputs(129)) and not (inputs(35));
    layer0_outputs(9478) <= not(inputs(74));
    layer0_outputs(9479) <= not(inputs(243)) or (inputs(255));
    layer0_outputs(9480) <= (inputs(102)) and not (inputs(144));
    layer0_outputs(9481) <= (inputs(129)) xor (inputs(131));
    layer0_outputs(9482) <= not(inputs(40)) or (inputs(174));
    layer0_outputs(9483) <= (inputs(30)) or (inputs(12));
    layer0_outputs(9484) <= not(inputs(122));
    layer0_outputs(9485) <= not((inputs(38)) xor (inputs(1)));
    layer0_outputs(9486) <= not(inputs(172)) or (inputs(150));
    layer0_outputs(9487) <= (inputs(41)) or (inputs(228));
    layer0_outputs(9488) <= not((inputs(193)) or (inputs(100)));
    layer0_outputs(9489) <= not((inputs(191)) or (inputs(194)));
    layer0_outputs(9490) <= inputs(101);
    layer0_outputs(9491) <= (inputs(76)) and (inputs(119));
    layer0_outputs(9492) <= not(inputs(151));
    layer0_outputs(9493) <= inputs(4);
    layer0_outputs(9494) <= '1';
    layer0_outputs(9495) <= (inputs(220)) or (inputs(212));
    layer0_outputs(9496) <= not((inputs(55)) and (inputs(52)));
    layer0_outputs(9497) <= not((inputs(211)) xor (inputs(106)));
    layer0_outputs(9498) <= (inputs(127)) or (inputs(2));
    layer0_outputs(9499) <= (inputs(151)) or (inputs(239));
    layer0_outputs(9500) <= not(inputs(18)) or (inputs(158));
    layer0_outputs(9501) <= (inputs(174)) xor (inputs(119));
    layer0_outputs(9502) <= not((inputs(32)) or (inputs(63)));
    layer0_outputs(9503) <= not(inputs(197)) or (inputs(172));
    layer0_outputs(9504) <= '1';
    layer0_outputs(9505) <= (inputs(135)) and not (inputs(144));
    layer0_outputs(9506) <= not((inputs(218)) or (inputs(82)));
    layer0_outputs(9507) <= not(inputs(161));
    layer0_outputs(9508) <= '0';
    layer0_outputs(9509) <= not(inputs(155));
    layer0_outputs(9510) <= inputs(46);
    layer0_outputs(9511) <= not(inputs(61));
    layer0_outputs(9512) <= (inputs(173)) xor (inputs(87));
    layer0_outputs(9513) <= not((inputs(208)) or (inputs(209)));
    layer0_outputs(9514) <= (inputs(75)) and not (inputs(71));
    layer0_outputs(9515) <= inputs(148);
    layer0_outputs(9516) <= not((inputs(247)) or (inputs(201)));
    layer0_outputs(9517) <= not(inputs(100));
    layer0_outputs(9518) <= not(inputs(130)) or (inputs(51));
    layer0_outputs(9519) <= not((inputs(129)) or (inputs(156)));
    layer0_outputs(9520) <= not((inputs(91)) or (inputs(96)));
    layer0_outputs(9521) <= not((inputs(66)) or (inputs(199)));
    layer0_outputs(9522) <= (inputs(225)) xor (inputs(196));
    layer0_outputs(9523) <= (inputs(117)) or (inputs(50));
    layer0_outputs(9524) <= (inputs(187)) and not (inputs(49));
    layer0_outputs(9525) <= not((inputs(234)) or (inputs(10)));
    layer0_outputs(9526) <= (inputs(234)) and not (inputs(59));
    layer0_outputs(9527) <= not((inputs(232)) xor (inputs(145)));
    layer0_outputs(9528) <= (inputs(238)) or (inputs(205));
    layer0_outputs(9529) <= (inputs(209)) or (inputs(25));
    layer0_outputs(9530) <= (inputs(213)) and not (inputs(112));
    layer0_outputs(9531) <= not((inputs(96)) xor (inputs(49)));
    layer0_outputs(9532) <= (inputs(205)) and (inputs(59));
    layer0_outputs(9533) <= not(inputs(92));
    layer0_outputs(9534) <= not(inputs(255));
    layer0_outputs(9535) <= not(inputs(53)) or (inputs(199));
    layer0_outputs(9536) <= (inputs(217)) and (inputs(92));
    layer0_outputs(9537) <= (inputs(21)) and not (inputs(68));
    layer0_outputs(9538) <= inputs(29);
    layer0_outputs(9539) <= not(inputs(239));
    layer0_outputs(9540) <= not(inputs(172));
    layer0_outputs(9541) <= not((inputs(160)) or (inputs(198)));
    layer0_outputs(9542) <= (inputs(132)) or (inputs(67));
    layer0_outputs(9543) <= (inputs(244)) and not (inputs(29));
    layer0_outputs(9544) <= not(inputs(168)) or (inputs(111));
    layer0_outputs(9545) <= not((inputs(105)) xor (inputs(177)));
    layer0_outputs(9546) <= not((inputs(178)) xor (inputs(1)));
    layer0_outputs(9547) <= (inputs(40)) and not (inputs(17));
    layer0_outputs(9548) <= not((inputs(11)) xor (inputs(44)));
    layer0_outputs(9549) <= (inputs(206)) or (inputs(186));
    layer0_outputs(9550) <= not((inputs(250)) or (inputs(147)));
    layer0_outputs(9551) <= (inputs(121)) or (inputs(31));
    layer0_outputs(9552) <= not((inputs(2)) or (inputs(232)));
    layer0_outputs(9553) <= (inputs(25)) xor (inputs(190));
    layer0_outputs(9554) <= inputs(56);
    layer0_outputs(9555) <= not((inputs(4)) or (inputs(123)));
    layer0_outputs(9556) <= not(inputs(77)) or (inputs(84));
    layer0_outputs(9557) <= not(inputs(134)) or (inputs(82));
    layer0_outputs(9558) <= (inputs(183)) or (inputs(117));
    layer0_outputs(9559) <= not(inputs(132)) or (inputs(0));
    layer0_outputs(9560) <= not(inputs(207));
    layer0_outputs(9561) <= not(inputs(195));
    layer0_outputs(9562) <= not((inputs(177)) or (inputs(156)));
    layer0_outputs(9563) <= (inputs(207)) or (inputs(2));
    layer0_outputs(9564) <= not(inputs(246));
    layer0_outputs(9565) <= not(inputs(184));
    layer0_outputs(9566) <= not((inputs(103)) xor (inputs(237)));
    layer0_outputs(9567) <= inputs(166);
    layer0_outputs(9568) <= inputs(72);
    layer0_outputs(9569) <= not(inputs(229));
    layer0_outputs(9570) <= (inputs(2)) and not (inputs(129));
    layer0_outputs(9571) <= not(inputs(147));
    layer0_outputs(9572) <= not(inputs(146));
    layer0_outputs(9573) <= '1';
    layer0_outputs(9574) <= not((inputs(163)) or (inputs(221)));
    layer0_outputs(9575) <= not(inputs(189));
    layer0_outputs(9576) <= (inputs(235)) and not (inputs(63));
    layer0_outputs(9577) <= not(inputs(189));
    layer0_outputs(9578) <= (inputs(154)) or (inputs(240));
    layer0_outputs(9579) <= not(inputs(116)) or (inputs(225));
    layer0_outputs(9580) <= not(inputs(112)) or (inputs(255));
    layer0_outputs(9581) <= not(inputs(55)) or (inputs(194));
    layer0_outputs(9582) <= inputs(182);
    layer0_outputs(9583) <= not((inputs(41)) and (inputs(177)));
    layer0_outputs(9584) <= not(inputs(10)) or (inputs(92));
    layer0_outputs(9585) <= not(inputs(104)) or (inputs(213));
    layer0_outputs(9586) <= inputs(230);
    layer0_outputs(9587) <= not(inputs(200));
    layer0_outputs(9588) <= not((inputs(115)) xor (inputs(86)));
    layer0_outputs(9589) <= not((inputs(53)) xor (inputs(70)));
    layer0_outputs(9590) <= not(inputs(46)) or (inputs(242));
    layer0_outputs(9591) <= (inputs(66)) and not (inputs(109));
    layer0_outputs(9592) <= (inputs(162)) and not (inputs(229));
    layer0_outputs(9593) <= (inputs(231)) or (inputs(194));
    layer0_outputs(9594) <= not((inputs(47)) or (inputs(99)));
    layer0_outputs(9595) <= (inputs(90)) xor (inputs(73));
    layer0_outputs(9596) <= not(inputs(110));
    layer0_outputs(9597) <= not(inputs(132));
    layer0_outputs(9598) <= not(inputs(58)) or (inputs(120));
    layer0_outputs(9599) <= inputs(121);
    layer0_outputs(9600) <= inputs(110);
    layer0_outputs(9601) <= not((inputs(74)) xor (inputs(43)));
    layer0_outputs(9602) <= not(inputs(132));
    layer0_outputs(9603) <= not(inputs(158));
    layer0_outputs(9604) <= inputs(32);
    layer0_outputs(9605) <= not(inputs(145)) or (inputs(28));
    layer0_outputs(9606) <= (inputs(224)) and (inputs(176));
    layer0_outputs(9607) <= (inputs(148)) and not (inputs(237));
    layer0_outputs(9608) <= not(inputs(246));
    layer0_outputs(9609) <= (inputs(95)) and (inputs(181));
    layer0_outputs(9610) <= not(inputs(145));
    layer0_outputs(9611) <= not(inputs(36)) or (inputs(176));
    layer0_outputs(9612) <= (inputs(48)) or (inputs(137));
    layer0_outputs(9613) <= not(inputs(206));
    layer0_outputs(9614) <= (inputs(173)) and (inputs(216));
    layer0_outputs(9615) <= (inputs(53)) and not (inputs(236));
    layer0_outputs(9616) <= inputs(218);
    layer0_outputs(9617) <= not(inputs(134)) or (inputs(173));
    layer0_outputs(9618) <= not((inputs(42)) or (inputs(72)));
    layer0_outputs(9619) <= not(inputs(143)) or (inputs(161));
    layer0_outputs(9620) <= inputs(208);
    layer0_outputs(9621) <= (inputs(241)) and not (inputs(142));
    layer0_outputs(9622) <= (inputs(251)) xor (inputs(249));
    layer0_outputs(9623) <= (inputs(123)) and not (inputs(216));
    layer0_outputs(9624) <= not((inputs(47)) or (inputs(136)));
    layer0_outputs(9625) <= inputs(131);
    layer0_outputs(9626) <= inputs(102);
    layer0_outputs(9627) <= not(inputs(213)) or (inputs(29));
    layer0_outputs(9628) <= (inputs(68)) and not (inputs(108));
    layer0_outputs(9629) <= (inputs(71)) and not (inputs(192));
    layer0_outputs(9630) <= not(inputs(97));
    layer0_outputs(9631) <= not((inputs(184)) xor (inputs(225)));
    layer0_outputs(9632) <= not(inputs(129)) or (inputs(13));
    layer0_outputs(9633) <= inputs(233);
    layer0_outputs(9634) <= not((inputs(91)) xor (inputs(137)));
    layer0_outputs(9635) <= not(inputs(187)) or (inputs(64));
    layer0_outputs(9636) <= (inputs(35)) xor (inputs(77));
    layer0_outputs(9637) <= not((inputs(156)) xor (inputs(16)));
    layer0_outputs(9638) <= not(inputs(136));
    layer0_outputs(9639) <= not(inputs(151));
    layer0_outputs(9640) <= not(inputs(157));
    layer0_outputs(9641) <= (inputs(12)) and not (inputs(154));
    layer0_outputs(9642) <= not((inputs(253)) or (inputs(196)));
    layer0_outputs(9643) <= not((inputs(130)) or (inputs(127)));
    layer0_outputs(9644) <= not(inputs(129));
    layer0_outputs(9645) <= not(inputs(158)) or (inputs(64));
    layer0_outputs(9646) <= (inputs(47)) or (inputs(13));
    layer0_outputs(9647) <= not(inputs(61));
    layer0_outputs(9648) <= not(inputs(235)) or (inputs(129));
    layer0_outputs(9649) <= (inputs(105)) or (inputs(8));
    layer0_outputs(9650) <= (inputs(133)) or (inputs(205));
    layer0_outputs(9651) <= (inputs(138)) xor (inputs(121));
    layer0_outputs(9652) <= (inputs(171)) xor (inputs(189));
    layer0_outputs(9653) <= inputs(120);
    layer0_outputs(9654) <= (inputs(131)) or (inputs(128));
    layer0_outputs(9655) <= not(inputs(183));
    layer0_outputs(9656) <= inputs(103);
    layer0_outputs(9657) <= (inputs(25)) xor (inputs(61));
    layer0_outputs(9658) <= not((inputs(23)) xor (inputs(210)));
    layer0_outputs(9659) <= (inputs(163)) or (inputs(26));
    layer0_outputs(9660) <= inputs(158);
    layer0_outputs(9661) <= (inputs(180)) and (inputs(239));
    layer0_outputs(9662) <= not((inputs(173)) or (inputs(144)));
    layer0_outputs(9663) <= not(inputs(151));
    layer0_outputs(9664) <= not(inputs(100));
    layer0_outputs(9665) <= (inputs(216)) and not (inputs(140));
    layer0_outputs(9666) <= (inputs(131)) and not (inputs(54));
    layer0_outputs(9667) <= (inputs(206)) or (inputs(52));
    layer0_outputs(9668) <= '0';
    layer0_outputs(9669) <= (inputs(171)) or (inputs(91));
    layer0_outputs(9670) <= (inputs(61)) xor (inputs(38));
    layer0_outputs(9671) <= not((inputs(1)) xor (inputs(46)));
    layer0_outputs(9672) <= not(inputs(98)) or (inputs(202));
    layer0_outputs(9673) <= inputs(157);
    layer0_outputs(9674) <= not((inputs(47)) and (inputs(15)));
    layer0_outputs(9675) <= not(inputs(176));
    layer0_outputs(9676) <= (inputs(31)) and not (inputs(137));
    layer0_outputs(9677) <= not(inputs(71)) or (inputs(154));
    layer0_outputs(9678) <= inputs(139);
    layer0_outputs(9679) <= not((inputs(107)) or (inputs(177)));
    layer0_outputs(9680) <= inputs(174);
    layer0_outputs(9681) <= '0';
    layer0_outputs(9682) <= not(inputs(73)) or (inputs(252));
    layer0_outputs(9683) <= (inputs(26)) xor (inputs(76));
    layer0_outputs(9684) <= not((inputs(202)) and (inputs(11)));
    layer0_outputs(9685) <= not((inputs(71)) or (inputs(164)));
    layer0_outputs(9686) <= (inputs(170)) and not (inputs(76));
    layer0_outputs(9687) <= inputs(220);
    layer0_outputs(9688) <= not(inputs(221));
    layer0_outputs(9689) <= not((inputs(5)) or (inputs(175)));
    layer0_outputs(9690) <= not(inputs(128)) or (inputs(3));
    layer0_outputs(9691) <= not((inputs(115)) and (inputs(23)));
    layer0_outputs(9692) <= (inputs(41)) and not (inputs(102));
    layer0_outputs(9693) <= inputs(93);
    layer0_outputs(9694) <= not(inputs(77));
    layer0_outputs(9695) <= (inputs(209)) or (inputs(165));
    layer0_outputs(9696) <= (inputs(135)) and (inputs(86));
    layer0_outputs(9697) <= not((inputs(32)) xor (inputs(99)));
    layer0_outputs(9698) <= not((inputs(233)) or (inputs(177)));
    layer0_outputs(9699) <= (inputs(105)) or (inputs(14));
    layer0_outputs(9700) <= '1';
    layer0_outputs(9701) <= inputs(111);
    layer0_outputs(9702) <= inputs(244);
    layer0_outputs(9703) <= (inputs(168)) or (inputs(86));
    layer0_outputs(9704) <= (inputs(252)) and not (inputs(93));
    layer0_outputs(9705) <= not(inputs(59));
    layer0_outputs(9706) <= not(inputs(28)) or (inputs(223));
    layer0_outputs(9707) <= inputs(8);
    layer0_outputs(9708) <= (inputs(69)) xor (inputs(66));
    layer0_outputs(9709) <= (inputs(81)) and (inputs(9));
    layer0_outputs(9710) <= inputs(70);
    layer0_outputs(9711) <= '0';
    layer0_outputs(9712) <= not(inputs(58));
    layer0_outputs(9713) <= inputs(213);
    layer0_outputs(9714) <= (inputs(4)) or (inputs(246));
    layer0_outputs(9715) <= not((inputs(235)) and (inputs(233)));
    layer0_outputs(9716) <= '1';
    layer0_outputs(9717) <= (inputs(143)) or (inputs(229));
    layer0_outputs(9718) <= not(inputs(49)) or (inputs(197));
    layer0_outputs(9719) <= inputs(245);
    layer0_outputs(9720) <= inputs(138);
    layer0_outputs(9721) <= not(inputs(1));
    layer0_outputs(9722) <= (inputs(230)) and not (inputs(237));
    layer0_outputs(9723) <= (inputs(246)) and not (inputs(165));
    layer0_outputs(9724) <= (inputs(176)) xor (inputs(67));
    layer0_outputs(9725) <= not(inputs(39)) or (inputs(59));
    layer0_outputs(9726) <= not(inputs(195));
    layer0_outputs(9727) <= '1';
    layer0_outputs(9728) <= not((inputs(136)) xor (inputs(222)));
    layer0_outputs(9729) <= not((inputs(14)) and (inputs(19)));
    layer0_outputs(9730) <= not(inputs(56)) or (inputs(147));
    layer0_outputs(9731) <= not((inputs(2)) or (inputs(73)));
    layer0_outputs(9732) <= (inputs(120)) and not (inputs(236));
    layer0_outputs(9733) <= not(inputs(153));
    layer0_outputs(9734) <= inputs(167);
    layer0_outputs(9735) <= (inputs(208)) or (inputs(96));
    layer0_outputs(9736) <= (inputs(20)) and not (inputs(223));
    layer0_outputs(9737) <= inputs(184);
    layer0_outputs(9738) <= not(inputs(21));
    layer0_outputs(9739) <= (inputs(103)) and not (inputs(224));
    layer0_outputs(9740) <= not(inputs(87)) or (inputs(35));
    layer0_outputs(9741) <= not((inputs(251)) or (inputs(173)));
    layer0_outputs(9742) <= inputs(73);
    layer0_outputs(9743) <= not((inputs(132)) xor (inputs(109)));
    layer0_outputs(9744) <= not(inputs(17)) or (inputs(227));
    layer0_outputs(9745) <= inputs(120);
    layer0_outputs(9746) <= (inputs(234)) and not (inputs(14));
    layer0_outputs(9747) <= not((inputs(150)) or (inputs(235)));
    layer0_outputs(9748) <= not((inputs(95)) or (inputs(75)));
    layer0_outputs(9749) <= (inputs(164)) or (inputs(51));
    layer0_outputs(9750) <= inputs(173);
    layer0_outputs(9751) <= not((inputs(74)) xor (inputs(47)));
    layer0_outputs(9752) <= (inputs(21)) xor (inputs(64));
    layer0_outputs(9753) <= (inputs(124)) and (inputs(20));
    layer0_outputs(9754) <= (inputs(44)) xor (inputs(40));
    layer0_outputs(9755) <= not(inputs(83));
    layer0_outputs(9756) <= not((inputs(126)) xor (inputs(71)));
    layer0_outputs(9757) <= (inputs(87)) or (inputs(218));
    layer0_outputs(9758) <= (inputs(99)) and not (inputs(254));
    layer0_outputs(9759) <= not(inputs(101));
    layer0_outputs(9760) <= (inputs(165)) or (inputs(108));
    layer0_outputs(9761) <= not(inputs(7)) or (inputs(176));
    layer0_outputs(9762) <= not((inputs(139)) or (inputs(84)));
    layer0_outputs(9763) <= (inputs(131)) and (inputs(122));
    layer0_outputs(9764) <= inputs(144);
    layer0_outputs(9765) <= not(inputs(102));
    layer0_outputs(9766) <= inputs(109);
    layer0_outputs(9767) <= (inputs(176)) and not (inputs(205));
    layer0_outputs(9768) <= inputs(26);
    layer0_outputs(9769) <= not((inputs(62)) or (inputs(34)));
    layer0_outputs(9770) <= not(inputs(40));
    layer0_outputs(9771) <= not(inputs(36));
    layer0_outputs(9772) <= inputs(249);
    layer0_outputs(9773) <= (inputs(107)) and not (inputs(67));
    layer0_outputs(9774) <= (inputs(98)) xor (inputs(171));
    layer0_outputs(9775) <= not(inputs(46));
    layer0_outputs(9776) <= not(inputs(46)) or (inputs(150));
    layer0_outputs(9777) <= not(inputs(131));
    layer0_outputs(9778) <= not(inputs(28)) or (inputs(15));
    layer0_outputs(9779) <= (inputs(185)) and not (inputs(2));
    layer0_outputs(9780) <= (inputs(248)) or (inputs(240));
    layer0_outputs(9781) <= not(inputs(199));
    layer0_outputs(9782) <= not(inputs(218));
    layer0_outputs(9783) <= (inputs(146)) or (inputs(85));
    layer0_outputs(9784) <= '0';
    layer0_outputs(9785) <= not((inputs(150)) and (inputs(37)));
    layer0_outputs(9786) <= (inputs(64)) or (inputs(39));
    layer0_outputs(9787) <= (inputs(35)) and (inputs(55));
    layer0_outputs(9788) <= not(inputs(117)) or (inputs(205));
    layer0_outputs(9789) <= not(inputs(25));
    layer0_outputs(9790) <= not((inputs(4)) xor (inputs(53)));
    layer0_outputs(9791) <= not((inputs(194)) or (inputs(216)));
    layer0_outputs(9792) <= (inputs(177)) xor (inputs(32));
    layer0_outputs(9793) <= not(inputs(159));
    layer0_outputs(9794) <= not(inputs(244)) or (inputs(119));
    layer0_outputs(9795) <= not(inputs(150)) or (inputs(12));
    layer0_outputs(9796) <= (inputs(23)) and not (inputs(163));
    layer0_outputs(9797) <= (inputs(218)) or (inputs(96));
    layer0_outputs(9798) <= (inputs(132)) xor (inputs(173));
    layer0_outputs(9799) <= inputs(198);
    layer0_outputs(9800) <= (inputs(70)) xor (inputs(49));
    layer0_outputs(9801) <= not(inputs(210));
    layer0_outputs(9802) <= (inputs(15)) or (inputs(55));
    layer0_outputs(9803) <= '0';
    layer0_outputs(9804) <= not((inputs(2)) or (inputs(89)));
    layer0_outputs(9805) <= not(inputs(158));
    layer0_outputs(9806) <= not(inputs(213)) or (inputs(33));
    layer0_outputs(9807) <= not(inputs(198)) or (inputs(44));
    layer0_outputs(9808) <= not((inputs(22)) or (inputs(246)));
    layer0_outputs(9809) <= not(inputs(94)) or (inputs(170));
    layer0_outputs(9810) <= (inputs(64)) or (inputs(5));
    layer0_outputs(9811) <= inputs(14);
    layer0_outputs(9812) <= (inputs(34)) xor (inputs(4));
    layer0_outputs(9813) <= not(inputs(81)) or (inputs(149));
    layer0_outputs(9814) <= not((inputs(207)) or (inputs(189)));
    layer0_outputs(9815) <= not(inputs(232)) or (inputs(88));
    layer0_outputs(9816) <= not(inputs(27));
    layer0_outputs(9817) <= inputs(252);
    layer0_outputs(9818) <= not(inputs(214));
    layer0_outputs(9819) <= not(inputs(152)) or (inputs(190));
    layer0_outputs(9820) <= (inputs(69)) and (inputs(187));
    layer0_outputs(9821) <= (inputs(244)) or (inputs(188));
    layer0_outputs(9822) <= not((inputs(209)) or (inputs(129)));
    layer0_outputs(9823) <= (inputs(99)) xor (inputs(145));
    layer0_outputs(9824) <= not(inputs(37)) or (inputs(166));
    layer0_outputs(9825) <= (inputs(60)) or (inputs(164));
    layer0_outputs(9826) <= not(inputs(41)) or (inputs(185));
    layer0_outputs(9827) <= not((inputs(89)) and (inputs(83)));
    layer0_outputs(9828) <= inputs(213);
    layer0_outputs(9829) <= inputs(182);
    layer0_outputs(9830) <= inputs(243);
    layer0_outputs(9831) <= not(inputs(65));
    layer0_outputs(9832) <= not(inputs(232)) or (inputs(103));
    layer0_outputs(9833) <= not((inputs(245)) or (inputs(6)));
    layer0_outputs(9834) <= (inputs(163)) or (inputs(26));
    layer0_outputs(9835) <= not(inputs(194)) or (inputs(30));
    layer0_outputs(9836) <= inputs(4);
    layer0_outputs(9837) <= inputs(148);
    layer0_outputs(9838) <= (inputs(219)) and (inputs(10));
    layer0_outputs(9839) <= inputs(202);
    layer0_outputs(9840) <= not(inputs(52)) or (inputs(61));
    layer0_outputs(9841) <= inputs(168);
    layer0_outputs(9842) <= not(inputs(196)) or (inputs(12));
    layer0_outputs(9843) <= not((inputs(92)) or (inputs(61)));
    layer0_outputs(9844) <= not(inputs(83));
    layer0_outputs(9845) <= inputs(84);
    layer0_outputs(9846) <= inputs(121);
    layer0_outputs(9847) <= inputs(234);
    layer0_outputs(9848) <= inputs(225);
    layer0_outputs(9849) <= not(inputs(27));
    layer0_outputs(9850) <= not((inputs(85)) xor (inputs(114)));
    layer0_outputs(9851) <= (inputs(17)) and not (inputs(74));
    layer0_outputs(9852) <= inputs(157);
    layer0_outputs(9853) <= inputs(48);
    layer0_outputs(9854) <= not(inputs(9)) or (inputs(2));
    layer0_outputs(9855) <= (inputs(58)) and not (inputs(66));
    layer0_outputs(9856) <= inputs(22);
    layer0_outputs(9857) <= inputs(219);
    layer0_outputs(9858) <= (inputs(46)) and not (inputs(167));
    layer0_outputs(9859) <= not((inputs(182)) and (inputs(123)));
    layer0_outputs(9860) <= not(inputs(30));
    layer0_outputs(9861) <= not(inputs(70)) or (inputs(252));
    layer0_outputs(9862) <= not(inputs(174)) or (inputs(103));
    layer0_outputs(9863) <= (inputs(146)) and not (inputs(34));
    layer0_outputs(9864) <= not(inputs(159));
    layer0_outputs(9865) <= (inputs(23)) or (inputs(136));
    layer0_outputs(9866) <= inputs(185);
    layer0_outputs(9867) <= not((inputs(159)) or (inputs(83)));
    layer0_outputs(9868) <= inputs(93);
    layer0_outputs(9869) <= not((inputs(172)) or (inputs(161)));
    layer0_outputs(9870) <= (inputs(112)) or (inputs(42));
    layer0_outputs(9871) <= (inputs(123)) or (inputs(129));
    layer0_outputs(9872) <= (inputs(159)) xor (inputs(216));
    layer0_outputs(9873) <= (inputs(49)) xor (inputs(100));
    layer0_outputs(9874) <= not(inputs(6));
    layer0_outputs(9875) <= '0';
    layer0_outputs(9876) <= inputs(33);
    layer0_outputs(9877) <= not(inputs(243)) or (inputs(54));
    layer0_outputs(9878) <= not(inputs(35));
    layer0_outputs(9879) <= inputs(218);
    layer0_outputs(9880) <= (inputs(195)) and not (inputs(105));
    layer0_outputs(9881) <= (inputs(19)) and not (inputs(242));
    layer0_outputs(9882) <= inputs(217);
    layer0_outputs(9883) <= not((inputs(250)) or (inputs(34)));
    layer0_outputs(9884) <= (inputs(48)) and not (inputs(154));
    layer0_outputs(9885) <= (inputs(130)) or (inputs(9));
    layer0_outputs(9886) <= (inputs(190)) or (inputs(111));
    layer0_outputs(9887) <= not(inputs(27));
    layer0_outputs(9888) <= not((inputs(168)) xor (inputs(253)));
    layer0_outputs(9889) <= not(inputs(68));
    layer0_outputs(9890) <= '0';
    layer0_outputs(9891) <= not((inputs(119)) or (inputs(120)));
    layer0_outputs(9892) <= not(inputs(114));
    layer0_outputs(9893) <= inputs(148);
    layer0_outputs(9894) <= inputs(247);
    layer0_outputs(9895) <= not(inputs(63));
    layer0_outputs(9896) <= (inputs(35)) and not (inputs(63));
    layer0_outputs(9897) <= (inputs(246)) and not (inputs(238));
    layer0_outputs(9898) <= inputs(19);
    layer0_outputs(9899) <= not(inputs(189));
    layer0_outputs(9900) <= not(inputs(129));
    layer0_outputs(9901) <= not(inputs(130));
    layer0_outputs(9902) <= not(inputs(167)) or (inputs(29));
    layer0_outputs(9903) <= (inputs(73)) or (inputs(139));
    layer0_outputs(9904) <= (inputs(173)) xor (inputs(108));
    layer0_outputs(9905) <= not(inputs(186)) or (inputs(31));
    layer0_outputs(9906) <= not(inputs(8));
    layer0_outputs(9907) <= (inputs(183)) or (inputs(99));
    layer0_outputs(9908) <= (inputs(209)) xor (inputs(166));
    layer0_outputs(9909) <= (inputs(209)) xor (inputs(80));
    layer0_outputs(9910) <= (inputs(160)) and (inputs(154));
    layer0_outputs(9911) <= not(inputs(8)) or (inputs(69));
    layer0_outputs(9912) <= inputs(235);
    layer0_outputs(9913) <= not(inputs(92));
    layer0_outputs(9914) <= '1';
    layer0_outputs(9915) <= not(inputs(120));
    layer0_outputs(9916) <= (inputs(149)) or (inputs(146));
    layer0_outputs(9917) <= '0';
    layer0_outputs(9918) <= not(inputs(53));
    layer0_outputs(9919) <= not(inputs(56));
    layer0_outputs(9920) <= inputs(68);
    layer0_outputs(9921) <= not(inputs(98));
    layer0_outputs(9922) <= (inputs(24)) and not (inputs(215));
    layer0_outputs(9923) <= (inputs(152)) and (inputs(94));
    layer0_outputs(9924) <= not(inputs(77));
    layer0_outputs(9925) <= (inputs(59)) and not (inputs(186));
    layer0_outputs(9926) <= (inputs(86)) or (inputs(93));
    layer0_outputs(9927) <= (inputs(26)) and not (inputs(176));
    layer0_outputs(9928) <= (inputs(196)) xor (inputs(104));
    layer0_outputs(9929) <= (inputs(85)) and not (inputs(234));
    layer0_outputs(9930) <= inputs(206);
    layer0_outputs(9931) <= (inputs(16)) and (inputs(125));
    layer0_outputs(9932) <= inputs(204);
    layer0_outputs(9933) <= not(inputs(202));
    layer0_outputs(9934) <= '0';
    layer0_outputs(9935) <= (inputs(85)) and not (inputs(214));
    layer0_outputs(9936) <= not(inputs(104)) or (inputs(81));
    layer0_outputs(9937) <= inputs(215);
    layer0_outputs(9938) <= not(inputs(201)) or (inputs(64));
    layer0_outputs(9939) <= not(inputs(86));
    layer0_outputs(9940) <= (inputs(65)) and not (inputs(175));
    layer0_outputs(9941) <= inputs(182);
    layer0_outputs(9942) <= not((inputs(27)) and (inputs(222)));
    layer0_outputs(9943) <= not(inputs(136)) or (inputs(222));
    layer0_outputs(9944) <= (inputs(136)) or (inputs(135));
    layer0_outputs(9945) <= (inputs(189)) xor (inputs(139));
    layer0_outputs(9946) <= not((inputs(101)) or (inputs(171)));
    layer0_outputs(9947) <= not((inputs(255)) xor (inputs(72)));
    layer0_outputs(9948) <= not(inputs(38)) or (inputs(250));
    layer0_outputs(9949) <= (inputs(182)) or (inputs(183));
    layer0_outputs(9950) <= (inputs(150)) or (inputs(167));
    layer0_outputs(9951) <= (inputs(208)) xor (inputs(152));
    layer0_outputs(9952) <= not(inputs(28)) or (inputs(236));
    layer0_outputs(9953) <= (inputs(16)) xor (inputs(6));
    layer0_outputs(9954) <= not(inputs(251)) or (inputs(160));
    layer0_outputs(9955) <= (inputs(184)) and not (inputs(53));
    layer0_outputs(9956) <= (inputs(68)) xor (inputs(36));
    layer0_outputs(9957) <= inputs(191);
    layer0_outputs(9958) <= (inputs(207)) xor (inputs(4));
    layer0_outputs(9959) <= not((inputs(95)) or (inputs(33)));
    layer0_outputs(9960) <= inputs(170);
    layer0_outputs(9961) <= (inputs(211)) and not (inputs(237));
    layer0_outputs(9962) <= not(inputs(149));
    layer0_outputs(9963) <= inputs(151);
    layer0_outputs(9964) <= not((inputs(52)) xor (inputs(251)));
    layer0_outputs(9965) <= not(inputs(202)) or (inputs(253));
    layer0_outputs(9966) <= not(inputs(137));
    layer0_outputs(9967) <= inputs(181);
    layer0_outputs(9968) <= (inputs(193)) or (inputs(221));
    layer0_outputs(9969) <= inputs(115);
    layer0_outputs(9970) <= (inputs(50)) or (inputs(107));
    layer0_outputs(9971) <= not(inputs(238));
    layer0_outputs(9972) <= not(inputs(26));
    layer0_outputs(9973) <= not((inputs(212)) and (inputs(209)));
    layer0_outputs(9974) <= not(inputs(141));
    layer0_outputs(9975) <= (inputs(198)) xor (inputs(180));
    layer0_outputs(9976) <= not((inputs(81)) xor (inputs(180)));
    layer0_outputs(9977) <= inputs(184);
    layer0_outputs(9978) <= (inputs(129)) xor (inputs(162));
    layer0_outputs(9979) <= (inputs(25)) xor (inputs(120));
    layer0_outputs(9980) <= inputs(140);
    layer0_outputs(9981) <= not(inputs(90));
    layer0_outputs(9982) <= not(inputs(133)) or (inputs(16));
    layer0_outputs(9983) <= inputs(174);
    layer0_outputs(9984) <= '0';
    layer0_outputs(9985) <= not((inputs(185)) xor (inputs(188)));
    layer0_outputs(9986) <= (inputs(46)) or (inputs(60));
    layer0_outputs(9987) <= not(inputs(79)) or (inputs(242));
    layer0_outputs(9988) <= (inputs(100)) and not (inputs(241));
    layer0_outputs(9989) <= not(inputs(98));
    layer0_outputs(9990) <= not(inputs(163));
    layer0_outputs(9991) <= inputs(109);
    layer0_outputs(9992) <= (inputs(119)) or (inputs(73));
    layer0_outputs(9993) <= not(inputs(53));
    layer0_outputs(9994) <= not((inputs(47)) or (inputs(34)));
    layer0_outputs(9995) <= (inputs(80)) xor (inputs(140));
    layer0_outputs(9996) <= not(inputs(145));
    layer0_outputs(9997) <= '1';
    layer0_outputs(9998) <= not(inputs(164));
    layer0_outputs(9999) <= not(inputs(246)) or (inputs(153));
    layer0_outputs(10000) <= '1';
    layer0_outputs(10001) <= (inputs(40)) and not (inputs(188));
    layer0_outputs(10002) <= not((inputs(215)) or (inputs(244)));
    layer0_outputs(10003) <= (inputs(144)) or (inputs(197));
    layer0_outputs(10004) <= inputs(168);
    layer0_outputs(10005) <= (inputs(51)) and not (inputs(240));
    layer0_outputs(10006) <= inputs(85);
    layer0_outputs(10007) <= not(inputs(32));
    layer0_outputs(10008) <= inputs(12);
    layer0_outputs(10009) <= inputs(181);
    layer0_outputs(10010) <= not(inputs(252));
    layer0_outputs(10011) <= (inputs(247)) and not (inputs(66));
    layer0_outputs(10012) <= not(inputs(42));
    layer0_outputs(10013) <= not(inputs(101)) or (inputs(254));
    layer0_outputs(10014) <= inputs(121);
    layer0_outputs(10015) <= inputs(52);
    layer0_outputs(10016) <= inputs(247);
    layer0_outputs(10017) <= inputs(19);
    layer0_outputs(10018) <= inputs(33);
    layer0_outputs(10019) <= inputs(90);
    layer0_outputs(10020) <= '1';
    layer0_outputs(10021) <= (inputs(35)) and not (inputs(237));
    layer0_outputs(10022) <= not(inputs(77));
    layer0_outputs(10023) <= not((inputs(101)) or (inputs(69)));
    layer0_outputs(10024) <= (inputs(226)) and (inputs(250));
    layer0_outputs(10025) <= inputs(249);
    layer0_outputs(10026) <= (inputs(17)) and not (inputs(183));
    layer0_outputs(10027) <= not((inputs(31)) or (inputs(177)));
    layer0_outputs(10028) <= not(inputs(180)) or (inputs(89));
    layer0_outputs(10029) <= (inputs(194)) or (inputs(195));
    layer0_outputs(10030) <= inputs(106);
    layer0_outputs(10031) <= not(inputs(85)) or (inputs(16));
    layer0_outputs(10032) <= not(inputs(182));
    layer0_outputs(10033) <= inputs(110);
    layer0_outputs(10034) <= not(inputs(207)) or (inputs(94));
    layer0_outputs(10035) <= inputs(35);
    layer0_outputs(10036) <= inputs(23);
    layer0_outputs(10037) <= (inputs(45)) and not (inputs(238));
    layer0_outputs(10038) <= not((inputs(168)) xor (inputs(104)));
    layer0_outputs(10039) <= (inputs(160)) xor (inputs(139));
    layer0_outputs(10040) <= (inputs(103)) or (inputs(178));
    layer0_outputs(10041) <= not((inputs(139)) and (inputs(139)));
    layer0_outputs(10042) <= inputs(23);
    layer0_outputs(10043) <= not(inputs(131));
    layer0_outputs(10044) <= not((inputs(34)) xor (inputs(244)));
    layer0_outputs(10045) <= (inputs(43)) and not (inputs(3));
    layer0_outputs(10046) <= not(inputs(95));
    layer0_outputs(10047) <= inputs(222);
    layer0_outputs(10048) <= inputs(37);
    layer0_outputs(10049) <= (inputs(231)) and (inputs(139));
    layer0_outputs(10050) <= '0';
    layer0_outputs(10051) <= not(inputs(66)) or (inputs(167));
    layer0_outputs(10052) <= (inputs(64)) xor (inputs(169));
    layer0_outputs(10053) <= not(inputs(173)) or (inputs(107));
    layer0_outputs(10054) <= (inputs(248)) and not (inputs(133));
    layer0_outputs(10055) <= not(inputs(224)) or (inputs(45));
    layer0_outputs(10056) <= not(inputs(90)) or (inputs(111));
    layer0_outputs(10057) <= (inputs(116)) or (inputs(51));
    layer0_outputs(10058) <= inputs(148);
    layer0_outputs(10059) <= (inputs(164)) and not (inputs(65));
    layer0_outputs(10060) <= not(inputs(148));
    layer0_outputs(10061) <= not(inputs(155)) or (inputs(153));
    layer0_outputs(10062) <= inputs(204);
    layer0_outputs(10063) <= inputs(200);
    layer0_outputs(10064) <= (inputs(200)) xor (inputs(232));
    layer0_outputs(10065) <= not(inputs(200));
    layer0_outputs(10066) <= not((inputs(25)) and (inputs(150)));
    layer0_outputs(10067) <= inputs(164);
    layer0_outputs(10068) <= (inputs(141)) xor (inputs(19));
    layer0_outputs(10069) <= not((inputs(142)) or (inputs(130)));
    layer0_outputs(10070) <= not(inputs(181)) or (inputs(253));
    layer0_outputs(10071) <= not(inputs(56)) or (inputs(233));
    layer0_outputs(10072) <= (inputs(25)) and not (inputs(149));
    layer0_outputs(10073) <= not(inputs(214));
    layer0_outputs(10074) <= (inputs(122)) and not (inputs(178));
    layer0_outputs(10075) <= inputs(161);
    layer0_outputs(10076) <= (inputs(170)) xor (inputs(162));
    layer0_outputs(10077) <= not(inputs(86));
    layer0_outputs(10078) <= not((inputs(13)) xor (inputs(223)));
    layer0_outputs(10079) <= (inputs(101)) and not (inputs(126));
    layer0_outputs(10080) <= inputs(120);
    layer0_outputs(10081) <= not(inputs(206)) or (inputs(69));
    layer0_outputs(10082) <= (inputs(133)) or (inputs(82));
    layer0_outputs(10083) <= inputs(131);
    layer0_outputs(10084) <= not((inputs(79)) or (inputs(71)));
    layer0_outputs(10085) <= inputs(114);
    layer0_outputs(10086) <= inputs(61);
    layer0_outputs(10087) <= (inputs(90)) and not (inputs(145));
    layer0_outputs(10088) <= (inputs(133)) or (inputs(238));
    layer0_outputs(10089) <= '1';
    layer0_outputs(10090) <= not(inputs(192)) or (inputs(221));
    layer0_outputs(10091) <= '0';
    layer0_outputs(10092) <= (inputs(236)) or (inputs(155));
    layer0_outputs(10093) <= not((inputs(127)) xor (inputs(247)));
    layer0_outputs(10094) <= (inputs(194)) and not (inputs(212));
    layer0_outputs(10095) <= '0';
    layer0_outputs(10096) <= not(inputs(109)) or (inputs(230));
    layer0_outputs(10097) <= not((inputs(190)) or (inputs(180)));
    layer0_outputs(10098) <= (inputs(112)) xor (inputs(44));
    layer0_outputs(10099) <= (inputs(167)) and not (inputs(129));
    layer0_outputs(10100) <= '0';
    layer0_outputs(10101) <= inputs(19);
    layer0_outputs(10102) <= (inputs(120)) and not (inputs(236));
    layer0_outputs(10103) <= (inputs(26)) and not (inputs(246));
    layer0_outputs(10104) <= inputs(114);
    layer0_outputs(10105) <= not((inputs(252)) or (inputs(233)));
    layer0_outputs(10106) <= not(inputs(247));
    layer0_outputs(10107) <= not(inputs(94));
    layer0_outputs(10108) <= not((inputs(22)) xor (inputs(82)));
    layer0_outputs(10109) <= not((inputs(35)) or (inputs(50)));
    layer0_outputs(10110) <= (inputs(14)) or (inputs(126));
    layer0_outputs(10111) <= (inputs(134)) and not (inputs(234));
    layer0_outputs(10112) <= (inputs(0)) and not (inputs(208));
    layer0_outputs(10113) <= not((inputs(230)) or (inputs(18)));
    layer0_outputs(10114) <= (inputs(122)) or (inputs(110));
    layer0_outputs(10115) <= not(inputs(99));
    layer0_outputs(10116) <= '1';
    layer0_outputs(10117) <= (inputs(100)) or (inputs(193));
    layer0_outputs(10118) <= not((inputs(239)) or (inputs(225)));
    layer0_outputs(10119) <= not((inputs(127)) or (inputs(43)));
    layer0_outputs(10120) <= inputs(114);
    layer0_outputs(10121) <= not((inputs(91)) xor (inputs(216)));
    layer0_outputs(10122) <= inputs(211);
    layer0_outputs(10123) <= not(inputs(232));
    layer0_outputs(10124) <= (inputs(127)) and not (inputs(115));
    layer0_outputs(10125) <= (inputs(149)) or (inputs(145));
    layer0_outputs(10126) <= not((inputs(205)) xor (inputs(104)));
    layer0_outputs(10127) <= (inputs(246)) or (inputs(2));
    layer0_outputs(10128) <= not((inputs(51)) or (inputs(195)));
    layer0_outputs(10129) <= (inputs(107)) and not (inputs(80));
    layer0_outputs(10130) <= (inputs(66)) or (inputs(195));
    layer0_outputs(10131) <= (inputs(184)) and not (inputs(61));
    layer0_outputs(10132) <= (inputs(246)) xor (inputs(4));
    layer0_outputs(10133) <= (inputs(163)) and not (inputs(78));
    layer0_outputs(10134) <= not(inputs(218));
    layer0_outputs(10135) <= (inputs(137)) and not (inputs(221));
    layer0_outputs(10136) <= not(inputs(215));
    layer0_outputs(10137) <= not(inputs(120));
    layer0_outputs(10138) <= (inputs(171)) and (inputs(48));
    layer0_outputs(10139) <= (inputs(239)) and not (inputs(161));
    layer0_outputs(10140) <= not((inputs(16)) and (inputs(198)));
    layer0_outputs(10141) <= not((inputs(226)) or (inputs(227)));
    layer0_outputs(10142) <= inputs(171);
    layer0_outputs(10143) <= (inputs(170)) or (inputs(59));
    layer0_outputs(10144) <= (inputs(86)) and not (inputs(152));
    layer0_outputs(10145) <= inputs(166);
    layer0_outputs(10146) <= not(inputs(153)) or (inputs(212));
    layer0_outputs(10147) <= not((inputs(221)) or (inputs(156)));
    layer0_outputs(10148) <= (inputs(103)) and (inputs(150));
    layer0_outputs(10149) <= inputs(89);
    layer0_outputs(10150) <= '0';
    layer0_outputs(10151) <= not((inputs(69)) or (inputs(99)));
    layer0_outputs(10152) <= (inputs(29)) or (inputs(154));
    layer0_outputs(10153) <= (inputs(234)) and not (inputs(240));
    layer0_outputs(10154) <= (inputs(182)) or (inputs(245));
    layer0_outputs(10155) <= not(inputs(106));
    layer0_outputs(10156) <= not(inputs(83)) or (inputs(109));
    layer0_outputs(10157) <= inputs(184);
    layer0_outputs(10158) <= not(inputs(140)) or (inputs(9));
    layer0_outputs(10159) <= (inputs(144)) and not (inputs(149));
    layer0_outputs(10160) <= not(inputs(211)) or (inputs(142));
    layer0_outputs(10161) <= not(inputs(122)) or (inputs(204));
    layer0_outputs(10162) <= not(inputs(3)) or (inputs(60));
    layer0_outputs(10163) <= (inputs(45)) and not (inputs(236));
    layer0_outputs(10164) <= inputs(214);
    layer0_outputs(10165) <= (inputs(30)) and not (inputs(177));
    layer0_outputs(10166) <= '0';
    layer0_outputs(10167) <= not((inputs(173)) or (inputs(163)));
    layer0_outputs(10168) <= not(inputs(155)) or (inputs(19));
    layer0_outputs(10169) <= '1';
    layer0_outputs(10170) <= (inputs(37)) or (inputs(81));
    layer0_outputs(10171) <= not(inputs(138)) or (inputs(244));
    layer0_outputs(10172) <= not((inputs(84)) xor (inputs(96)));
    layer0_outputs(10173) <= '0';
    layer0_outputs(10174) <= inputs(77);
    layer0_outputs(10175) <= (inputs(129)) xor (inputs(68));
    layer0_outputs(10176) <= (inputs(141)) or (inputs(220));
    layer0_outputs(10177) <= (inputs(139)) and not (inputs(95));
    layer0_outputs(10178) <= not((inputs(84)) or (inputs(202)));
    layer0_outputs(10179) <= not(inputs(167)) or (inputs(249));
    layer0_outputs(10180) <= not(inputs(184));
    layer0_outputs(10181) <= not(inputs(93)) or (inputs(96));
    layer0_outputs(10182) <= (inputs(4)) or (inputs(120));
    layer0_outputs(10183) <= not(inputs(131));
    layer0_outputs(10184) <= (inputs(177)) or (inputs(214));
    layer0_outputs(10185) <= not(inputs(15));
    layer0_outputs(10186) <= '1';
    layer0_outputs(10187) <= not((inputs(193)) and (inputs(67)));
    layer0_outputs(10188) <= (inputs(181)) or (inputs(227));
    layer0_outputs(10189) <= (inputs(19)) or (inputs(227));
    layer0_outputs(10190) <= not(inputs(99));
    layer0_outputs(10191) <= (inputs(86)) xor (inputs(161));
    layer0_outputs(10192) <= inputs(242);
    layer0_outputs(10193) <= not(inputs(78)) or (inputs(28));
    layer0_outputs(10194) <= not(inputs(217)) or (inputs(70));
    layer0_outputs(10195) <= (inputs(33)) or (inputs(48));
    layer0_outputs(10196) <= '1';
    layer0_outputs(10197) <= inputs(237);
    layer0_outputs(10198) <= not(inputs(2));
    layer0_outputs(10199) <= (inputs(189)) and not (inputs(44));
    layer0_outputs(10200) <= inputs(157);
    layer0_outputs(10201) <= (inputs(111)) or (inputs(2));
    layer0_outputs(10202) <= (inputs(115)) or (inputs(198));
    layer0_outputs(10203) <= not(inputs(122));
    layer0_outputs(10204) <= (inputs(135)) and (inputs(11));
    layer0_outputs(10205) <= (inputs(170)) or (inputs(105));
    layer0_outputs(10206) <= not((inputs(195)) xor (inputs(197)));
    layer0_outputs(10207) <= not(inputs(242));
    layer0_outputs(10208) <= (inputs(227)) and not (inputs(0));
    layer0_outputs(10209) <= not(inputs(126));
    layer0_outputs(10210) <= inputs(234);
    layer0_outputs(10211) <= not((inputs(177)) xor (inputs(113)));
    layer0_outputs(10212) <= '0';
    layer0_outputs(10213) <= not(inputs(210));
    layer0_outputs(10214) <= (inputs(232)) and not (inputs(45));
    layer0_outputs(10215) <= (inputs(19)) xor (inputs(103));
    layer0_outputs(10216) <= not((inputs(86)) or (inputs(200)));
    layer0_outputs(10217) <= inputs(183);
    layer0_outputs(10218) <= not((inputs(31)) or (inputs(123)));
    layer0_outputs(10219) <= not((inputs(147)) xor (inputs(18)));
    layer0_outputs(10220) <= (inputs(46)) and not (inputs(244));
    layer0_outputs(10221) <= not(inputs(144)) or (inputs(221));
    layer0_outputs(10222) <= (inputs(166)) and not (inputs(244));
    layer0_outputs(10223) <= not((inputs(188)) or (inputs(255)));
    layer0_outputs(10224) <= (inputs(113)) xor (inputs(100));
    layer0_outputs(10225) <= not((inputs(95)) or (inputs(208)));
    layer0_outputs(10226) <= not(inputs(245)) or (inputs(1));
    layer0_outputs(10227) <= '1';
    layer0_outputs(10228) <= not((inputs(70)) xor (inputs(201)));
    layer0_outputs(10229) <= (inputs(239)) xor (inputs(63));
    layer0_outputs(10230) <= not((inputs(169)) or (inputs(127)));
    layer0_outputs(10231) <= not((inputs(38)) or (inputs(35)));
    layer0_outputs(10232) <= inputs(144);
    layer0_outputs(10233) <= (inputs(192)) or (inputs(225));
    layer0_outputs(10234) <= not((inputs(25)) or (inputs(8)));
    layer0_outputs(10235) <= inputs(84);
    layer0_outputs(10236) <= (inputs(214)) and not (inputs(93));
    layer0_outputs(10237) <= (inputs(132)) and not (inputs(80));
    layer0_outputs(10238) <= (inputs(140)) and (inputs(0));
    layer0_outputs(10239) <= not(inputs(85));
    layer1_outputs(0) <= layer0_outputs(4139);
    layer1_outputs(1) <= not(layer0_outputs(2922)) or (layer0_outputs(1196));
    layer1_outputs(2) <= layer0_outputs(3858);
    layer1_outputs(3) <= not(layer0_outputs(4282));
    layer1_outputs(4) <= not(layer0_outputs(4140));
    layer1_outputs(5) <= layer0_outputs(5458);
    layer1_outputs(6) <= (layer0_outputs(6133)) or (layer0_outputs(8679));
    layer1_outputs(7) <= not((layer0_outputs(5693)) or (layer0_outputs(9335)));
    layer1_outputs(8) <= (layer0_outputs(4004)) and (layer0_outputs(9310));
    layer1_outputs(9) <= not(layer0_outputs(9215)) or (layer0_outputs(7883));
    layer1_outputs(10) <= not(layer0_outputs(2319)) or (layer0_outputs(8529));
    layer1_outputs(11) <= layer0_outputs(291);
    layer1_outputs(12) <= layer0_outputs(932);
    layer1_outputs(13) <= (layer0_outputs(239)) xor (layer0_outputs(3763));
    layer1_outputs(14) <= not(layer0_outputs(336)) or (layer0_outputs(7458));
    layer1_outputs(15) <= (layer0_outputs(2759)) and (layer0_outputs(3848));
    layer1_outputs(16) <= (layer0_outputs(2376)) xor (layer0_outputs(6504));
    layer1_outputs(17) <= (layer0_outputs(7012)) xor (layer0_outputs(5921));
    layer1_outputs(18) <= (layer0_outputs(7365)) and (layer0_outputs(5167));
    layer1_outputs(19) <= not(layer0_outputs(7718));
    layer1_outputs(20) <= (layer0_outputs(1034)) or (layer0_outputs(512));
    layer1_outputs(21) <= (layer0_outputs(8807)) and not (layer0_outputs(3104));
    layer1_outputs(22) <= not(layer0_outputs(5641));
    layer1_outputs(23) <= not((layer0_outputs(9576)) xor (layer0_outputs(6451)));
    layer1_outputs(24) <= (layer0_outputs(3279)) and not (layer0_outputs(3681));
    layer1_outputs(25) <= not(layer0_outputs(8212)) or (layer0_outputs(5199));
    layer1_outputs(26) <= layer0_outputs(10185);
    layer1_outputs(27) <= (layer0_outputs(72)) xor (layer0_outputs(1969));
    layer1_outputs(28) <= not((layer0_outputs(7519)) and (layer0_outputs(2612)));
    layer1_outputs(29) <= not((layer0_outputs(1863)) and (layer0_outputs(1834)));
    layer1_outputs(30) <= (layer0_outputs(7288)) and (layer0_outputs(2285));
    layer1_outputs(31) <= '0';
    layer1_outputs(32) <= (layer0_outputs(7733)) or (layer0_outputs(5266));
    layer1_outputs(33) <= not((layer0_outputs(10030)) xor (layer0_outputs(9720)));
    layer1_outputs(34) <= not(layer0_outputs(6682));
    layer1_outputs(35) <= (layer0_outputs(3703)) and not (layer0_outputs(5791));
    layer1_outputs(36) <= (layer0_outputs(3481)) xor (layer0_outputs(5184));
    layer1_outputs(37) <= not(layer0_outputs(7209)) or (layer0_outputs(4901));
    layer1_outputs(38) <= not(layer0_outputs(7080)) or (layer0_outputs(7792));
    layer1_outputs(39) <= not(layer0_outputs(1780));
    layer1_outputs(40) <= layer0_outputs(10205);
    layer1_outputs(41) <= (layer0_outputs(1332)) or (layer0_outputs(7489));
    layer1_outputs(42) <= (layer0_outputs(2735)) or (layer0_outputs(6512));
    layer1_outputs(43) <= not((layer0_outputs(5988)) and (layer0_outputs(3493)));
    layer1_outputs(44) <= not((layer0_outputs(9365)) xor (layer0_outputs(10170)));
    layer1_outputs(45) <= not((layer0_outputs(583)) and (layer0_outputs(9227)));
    layer1_outputs(46) <= not(layer0_outputs(8635)) or (layer0_outputs(6666));
    layer1_outputs(47) <= not(layer0_outputs(1161));
    layer1_outputs(48) <= not(layer0_outputs(4887));
    layer1_outputs(49) <= (layer0_outputs(965)) and not (layer0_outputs(1753));
    layer1_outputs(50) <= layer0_outputs(7082);
    layer1_outputs(51) <= (layer0_outputs(4738)) and not (layer0_outputs(3699));
    layer1_outputs(52) <= not((layer0_outputs(5834)) xor (layer0_outputs(4510)));
    layer1_outputs(53) <= not((layer0_outputs(3270)) xor (layer0_outputs(4028)));
    layer1_outputs(54) <= (layer0_outputs(4071)) and not (layer0_outputs(8469));
    layer1_outputs(55) <= (layer0_outputs(6529)) or (layer0_outputs(2041));
    layer1_outputs(56) <= layer0_outputs(1158);
    layer1_outputs(57) <= layer0_outputs(2525);
    layer1_outputs(58) <= layer0_outputs(6671);
    layer1_outputs(59) <= not(layer0_outputs(3075));
    layer1_outputs(60) <= (layer0_outputs(5159)) or (layer0_outputs(6439));
    layer1_outputs(61) <= not((layer0_outputs(953)) and (layer0_outputs(2938)));
    layer1_outputs(62) <= not(layer0_outputs(4461));
    layer1_outputs(63) <= (layer0_outputs(3468)) xor (layer0_outputs(8286));
    layer1_outputs(64) <= layer0_outputs(2659);
    layer1_outputs(65) <= layer0_outputs(902);
    layer1_outputs(66) <= not((layer0_outputs(3575)) or (layer0_outputs(1410)));
    layer1_outputs(67) <= layer0_outputs(8481);
    layer1_outputs(68) <= not((layer0_outputs(2883)) and (layer0_outputs(920)));
    layer1_outputs(69) <= (layer0_outputs(6595)) and not (layer0_outputs(6724));
    layer1_outputs(70) <= not(layer0_outputs(5789));
    layer1_outputs(71) <= not((layer0_outputs(33)) or (layer0_outputs(8845)));
    layer1_outputs(72) <= layer0_outputs(4413);
    layer1_outputs(73) <= not(layer0_outputs(3000));
    layer1_outputs(74) <= (layer0_outputs(3713)) xor (layer0_outputs(6406));
    layer1_outputs(75) <= layer0_outputs(8802);
    layer1_outputs(76) <= not(layer0_outputs(361));
    layer1_outputs(77) <= not(layer0_outputs(1101));
    layer1_outputs(78) <= (layer0_outputs(1988)) or (layer0_outputs(7245));
    layer1_outputs(79) <= not(layer0_outputs(8366));
    layer1_outputs(80) <= (layer0_outputs(1962)) or (layer0_outputs(486));
    layer1_outputs(81) <= not(layer0_outputs(43));
    layer1_outputs(82) <= not(layer0_outputs(2502));
    layer1_outputs(83) <= (layer0_outputs(6319)) or (layer0_outputs(2903));
    layer1_outputs(84) <= (layer0_outputs(4502)) or (layer0_outputs(8137));
    layer1_outputs(85) <= '0';
    layer1_outputs(86) <= layer0_outputs(715);
    layer1_outputs(87) <= (layer0_outputs(8697)) and (layer0_outputs(2668));
    layer1_outputs(88) <= not((layer0_outputs(8528)) or (layer0_outputs(7161)));
    layer1_outputs(89) <= (layer0_outputs(4621)) and not (layer0_outputs(486));
    layer1_outputs(90) <= not(layer0_outputs(2940)) or (layer0_outputs(661));
    layer1_outputs(91) <= not(layer0_outputs(6745)) or (layer0_outputs(9418));
    layer1_outputs(92) <= (layer0_outputs(4503)) and not (layer0_outputs(5053));
    layer1_outputs(93) <= layer0_outputs(8115);
    layer1_outputs(94) <= not(layer0_outputs(8832)) or (layer0_outputs(3994));
    layer1_outputs(95) <= layer0_outputs(1519);
    layer1_outputs(96) <= layer0_outputs(1697);
    layer1_outputs(97) <= not(layer0_outputs(5344)) or (layer0_outputs(4564));
    layer1_outputs(98) <= not(layer0_outputs(6559)) or (layer0_outputs(2381));
    layer1_outputs(99) <= (layer0_outputs(255)) and not (layer0_outputs(1993));
    layer1_outputs(100) <= layer0_outputs(3806);
    layer1_outputs(101) <= layer0_outputs(1860);
    layer1_outputs(102) <= '1';
    layer1_outputs(103) <= (layer0_outputs(6589)) and (layer0_outputs(1602));
    layer1_outputs(104) <= not(layer0_outputs(1877));
    layer1_outputs(105) <= (layer0_outputs(8294)) xor (layer0_outputs(8990));
    layer1_outputs(106) <= not((layer0_outputs(3523)) and (layer0_outputs(2616)));
    layer1_outputs(107) <= not((layer0_outputs(6831)) and (layer0_outputs(6939)));
    layer1_outputs(108) <= not((layer0_outputs(1509)) xor (layer0_outputs(2592)));
    layer1_outputs(109) <= not(layer0_outputs(4993)) or (layer0_outputs(8236));
    layer1_outputs(110) <= not((layer0_outputs(3490)) and (layer0_outputs(956)));
    layer1_outputs(111) <= not(layer0_outputs(7343));
    layer1_outputs(112) <= layer0_outputs(1151);
    layer1_outputs(113) <= (layer0_outputs(10057)) xor (layer0_outputs(5221));
    layer1_outputs(114) <= (layer0_outputs(2910)) and (layer0_outputs(7511));
    layer1_outputs(115) <= (layer0_outputs(6399)) xor (layer0_outputs(8524));
    layer1_outputs(116) <= not(layer0_outputs(3770));
    layer1_outputs(117) <= not((layer0_outputs(1246)) or (layer0_outputs(9746)));
    layer1_outputs(118) <= (layer0_outputs(3578)) and not (layer0_outputs(6582));
    layer1_outputs(119) <= (layer0_outputs(8907)) and (layer0_outputs(4447));
    layer1_outputs(120) <= (layer0_outputs(5572)) and (layer0_outputs(8933));
    layer1_outputs(121) <= not(layer0_outputs(3740));
    layer1_outputs(122) <= (layer0_outputs(7284)) or (layer0_outputs(6304));
    layer1_outputs(123) <= (layer0_outputs(4009)) or (layer0_outputs(1645));
    layer1_outputs(124) <= not(layer0_outputs(1893));
    layer1_outputs(125) <= not(layer0_outputs(3819));
    layer1_outputs(126) <= not(layer0_outputs(2030));
    layer1_outputs(127) <= not(layer0_outputs(8403)) or (layer0_outputs(9824));
    layer1_outputs(128) <= (layer0_outputs(7068)) and (layer0_outputs(3722));
    layer1_outputs(129) <= not(layer0_outputs(3672));
    layer1_outputs(130) <= layer0_outputs(8748);
    layer1_outputs(131) <= not((layer0_outputs(8112)) or (layer0_outputs(1455)));
    layer1_outputs(132) <= not(layer0_outputs(1434));
    layer1_outputs(133) <= (layer0_outputs(1034)) and not (layer0_outputs(2665));
    layer1_outputs(134) <= '1';
    layer1_outputs(135) <= layer0_outputs(4594);
    layer1_outputs(136) <= (layer0_outputs(8690)) and not (layer0_outputs(9519));
    layer1_outputs(137) <= (layer0_outputs(6139)) and not (layer0_outputs(10139));
    layer1_outputs(138) <= layer0_outputs(6045);
    layer1_outputs(139) <= (layer0_outputs(5437)) or (layer0_outputs(3438));
    layer1_outputs(140) <= not(layer0_outputs(3805));
    layer1_outputs(141) <= not(layer0_outputs(5093));
    layer1_outputs(142) <= not((layer0_outputs(7831)) xor (layer0_outputs(684)));
    layer1_outputs(143) <= (layer0_outputs(7191)) and not (layer0_outputs(4744));
    layer1_outputs(144) <= not(layer0_outputs(10128)) or (layer0_outputs(4248));
    layer1_outputs(145) <= not((layer0_outputs(6739)) or (layer0_outputs(6970)));
    layer1_outputs(146) <= (layer0_outputs(6803)) and (layer0_outputs(9861));
    layer1_outputs(147) <= (layer0_outputs(165)) xor (layer0_outputs(7791));
    layer1_outputs(148) <= not(layer0_outputs(5297));
    layer1_outputs(149) <= not(layer0_outputs(10031));
    layer1_outputs(150) <= (layer0_outputs(2264)) and not (layer0_outputs(9419));
    layer1_outputs(151) <= layer0_outputs(3162);
    layer1_outputs(152) <= (layer0_outputs(2849)) and not (layer0_outputs(6679));
    layer1_outputs(153) <= not(layer0_outputs(7171));
    layer1_outputs(154) <= layer0_outputs(9541);
    layer1_outputs(155) <= not(layer0_outputs(2993));
    layer1_outputs(156) <= (layer0_outputs(4529)) and not (layer0_outputs(5019));
    layer1_outputs(157) <= '1';
    layer1_outputs(158) <= not(layer0_outputs(3512));
    layer1_outputs(159) <= (layer0_outputs(7772)) xor (layer0_outputs(9680));
    layer1_outputs(160) <= not(layer0_outputs(5139));
    layer1_outputs(161) <= not(layer0_outputs(9478));
    layer1_outputs(162) <= not(layer0_outputs(4643));
    layer1_outputs(163) <= not(layer0_outputs(4111));
    layer1_outputs(164) <= (layer0_outputs(7846)) or (layer0_outputs(10142));
    layer1_outputs(165) <= (layer0_outputs(7297)) and not (layer0_outputs(8792));
    layer1_outputs(166) <= layer0_outputs(1135);
    layer1_outputs(167) <= layer0_outputs(6276);
    layer1_outputs(168) <= not(layer0_outputs(7026));
    layer1_outputs(169) <= layer0_outputs(3779);
    layer1_outputs(170) <= (layer0_outputs(2496)) or (layer0_outputs(9784));
    layer1_outputs(171) <= layer0_outputs(1292);
    layer1_outputs(172) <= not(layer0_outputs(5317));
    layer1_outputs(173) <= layer0_outputs(6032);
    layer1_outputs(174) <= not(layer0_outputs(9082));
    layer1_outputs(175) <= (layer0_outputs(3883)) and (layer0_outputs(9605));
    layer1_outputs(176) <= not(layer0_outputs(7498));
    layer1_outputs(177) <= (layer0_outputs(7565)) and (layer0_outputs(860));
    layer1_outputs(178) <= (layer0_outputs(4970)) and not (layer0_outputs(3242));
    layer1_outputs(179) <= (layer0_outputs(9307)) and not (layer0_outputs(2137));
    layer1_outputs(180) <= not(layer0_outputs(9734));
    layer1_outputs(181) <= not(layer0_outputs(4693));
    layer1_outputs(182) <= (layer0_outputs(4527)) and (layer0_outputs(9318));
    layer1_outputs(183) <= (layer0_outputs(500)) or (layer0_outputs(7281));
    layer1_outputs(184) <= not((layer0_outputs(3361)) or (layer0_outputs(1501)));
    layer1_outputs(185) <= layer0_outputs(1688);
    layer1_outputs(186) <= layer0_outputs(4553);
    layer1_outputs(187) <= (layer0_outputs(2263)) and not (layer0_outputs(1844));
    layer1_outputs(188) <= not((layer0_outputs(1767)) or (layer0_outputs(2600)));
    layer1_outputs(189) <= not((layer0_outputs(1215)) and (layer0_outputs(4598)));
    layer1_outputs(190) <= (layer0_outputs(8454)) and (layer0_outputs(9371));
    layer1_outputs(191) <= layer0_outputs(3928);
    layer1_outputs(192) <= layer0_outputs(6913);
    layer1_outputs(193) <= not(layer0_outputs(2382)) or (layer0_outputs(2598));
    layer1_outputs(194) <= (layer0_outputs(8800)) and not (layer0_outputs(8209));
    layer1_outputs(195) <= not((layer0_outputs(5338)) xor (layer0_outputs(2571)));
    layer1_outputs(196) <= not(layer0_outputs(2797)) or (layer0_outputs(2155));
    layer1_outputs(197) <= (layer0_outputs(9417)) or (layer0_outputs(2856));
    layer1_outputs(198) <= layer0_outputs(7003);
    layer1_outputs(199) <= not(layer0_outputs(9588));
    layer1_outputs(200) <= (layer0_outputs(9802)) xor (layer0_outputs(1646));
    layer1_outputs(201) <= layer0_outputs(7433);
    layer1_outputs(202) <= not(layer0_outputs(6674));
    layer1_outputs(203) <= not(layer0_outputs(9843));
    layer1_outputs(204) <= layer0_outputs(3103);
    layer1_outputs(205) <= not(layer0_outputs(8370)) or (layer0_outputs(7113));
    layer1_outputs(206) <= (layer0_outputs(469)) and not (layer0_outputs(5540));
    layer1_outputs(207) <= layer0_outputs(9389);
    layer1_outputs(208) <= layer0_outputs(914);
    layer1_outputs(209) <= layer0_outputs(9967);
    layer1_outputs(210) <= (layer0_outputs(8842)) or (layer0_outputs(9980));
    layer1_outputs(211) <= not(layer0_outputs(5737));
    layer1_outputs(212) <= not(layer0_outputs(4453)) or (layer0_outputs(3967));
    layer1_outputs(213) <= (layer0_outputs(5644)) and not (layer0_outputs(6668));
    layer1_outputs(214) <= (layer0_outputs(8173)) and not (layer0_outputs(4540));
    layer1_outputs(215) <= (layer0_outputs(10222)) or (layer0_outputs(4638));
    layer1_outputs(216) <= not(layer0_outputs(1570)) or (layer0_outputs(1156));
    layer1_outputs(217) <= not((layer0_outputs(6423)) or (layer0_outputs(8923)));
    layer1_outputs(218) <= not(layer0_outputs(3678));
    layer1_outputs(219) <= (layer0_outputs(8944)) and (layer0_outputs(1206));
    layer1_outputs(220) <= not(layer0_outputs(5315)) or (layer0_outputs(3785));
    layer1_outputs(221) <= (layer0_outputs(9378)) or (layer0_outputs(6384));
    layer1_outputs(222) <= (layer0_outputs(210)) and not (layer0_outputs(8699));
    layer1_outputs(223) <= (layer0_outputs(9302)) or (layer0_outputs(5494));
    layer1_outputs(224) <= not((layer0_outputs(563)) or (layer0_outputs(5377)));
    layer1_outputs(225) <= (layer0_outputs(5263)) xor (layer0_outputs(7155));
    layer1_outputs(226) <= not(layer0_outputs(1882));
    layer1_outputs(227) <= not((layer0_outputs(5498)) or (layer0_outputs(5947)));
    layer1_outputs(228) <= (layer0_outputs(4958)) and (layer0_outputs(9398));
    layer1_outputs(229) <= (layer0_outputs(3926)) or (layer0_outputs(6392));
    layer1_outputs(230) <= (layer0_outputs(767)) and not (layer0_outputs(9762));
    layer1_outputs(231) <= layer0_outputs(4571);
    layer1_outputs(232) <= not(layer0_outputs(5564));
    layer1_outputs(233) <= (layer0_outputs(10161)) and not (layer0_outputs(871));
    layer1_outputs(234) <= not((layer0_outputs(1493)) and (layer0_outputs(2678)));
    layer1_outputs(235) <= not(layer0_outputs(1505));
    layer1_outputs(236) <= layer0_outputs(7766);
    layer1_outputs(237) <= (layer0_outputs(9751)) and not (layer0_outputs(2708));
    layer1_outputs(238) <= not(layer0_outputs(9235));
    layer1_outputs(239) <= not(layer0_outputs(6939));
    layer1_outputs(240) <= not((layer0_outputs(1549)) xor (layer0_outputs(5161)));
    layer1_outputs(241) <= not(layer0_outputs(1085));
    layer1_outputs(242) <= not(layer0_outputs(800)) or (layer0_outputs(8378));
    layer1_outputs(243) <= layer0_outputs(8420);
    layer1_outputs(244) <= not(layer0_outputs(4682)) or (layer0_outputs(4957));
    layer1_outputs(245) <= not(layer0_outputs(1599));
    layer1_outputs(246) <= (layer0_outputs(9670)) xor (layer0_outputs(2769));
    layer1_outputs(247) <= not((layer0_outputs(3567)) or (layer0_outputs(8184)));
    layer1_outputs(248) <= not((layer0_outputs(6184)) xor (layer0_outputs(1024)));
    layer1_outputs(249) <= (layer0_outputs(1319)) and not (layer0_outputs(2857));
    layer1_outputs(250) <= not((layer0_outputs(34)) xor (layer0_outputs(5867)));
    layer1_outputs(251) <= not((layer0_outputs(9625)) or (layer0_outputs(6357)));
    layer1_outputs(252) <= (layer0_outputs(3172)) and not (layer0_outputs(7743));
    layer1_outputs(253) <= (layer0_outputs(5738)) and (layer0_outputs(592));
    layer1_outputs(254) <= layer0_outputs(2402);
    layer1_outputs(255) <= (layer0_outputs(6909)) or (layer0_outputs(97));
    layer1_outputs(256) <= (layer0_outputs(6514)) and (layer0_outputs(3673));
    layer1_outputs(257) <= not((layer0_outputs(7322)) and (layer0_outputs(4807)));
    layer1_outputs(258) <= (layer0_outputs(5884)) or (layer0_outputs(9412));
    layer1_outputs(259) <= layer0_outputs(1909);
    layer1_outputs(260) <= not(layer0_outputs(9996));
    layer1_outputs(261) <= not(layer0_outputs(6686)) or (layer0_outputs(583));
    layer1_outputs(262) <= not(layer0_outputs(8996));
    layer1_outputs(263) <= layer0_outputs(6122);
    layer1_outputs(264) <= (layer0_outputs(9186)) and not (layer0_outputs(2613));
    layer1_outputs(265) <= not(layer0_outputs(217));
    layer1_outputs(266) <= layer0_outputs(9682);
    layer1_outputs(267) <= layer0_outputs(5474);
    layer1_outputs(268) <= '1';
    layer1_outputs(269) <= (layer0_outputs(3884)) or (layer0_outputs(7825));
    layer1_outputs(270) <= layer0_outputs(2892);
    layer1_outputs(271) <= not(layer0_outputs(1449)) or (layer0_outputs(9301));
    layer1_outputs(272) <= not(layer0_outputs(9277)) or (layer0_outputs(716));
    layer1_outputs(273) <= (layer0_outputs(3121)) xor (layer0_outputs(5243));
    layer1_outputs(274) <= layer0_outputs(6800);
    layer1_outputs(275) <= (layer0_outputs(5715)) and not (layer0_outputs(3627));
    layer1_outputs(276) <= not(layer0_outputs(127));
    layer1_outputs(277) <= (layer0_outputs(3627)) or (layer0_outputs(7768));
    layer1_outputs(278) <= (layer0_outputs(7900)) and not (layer0_outputs(2811));
    layer1_outputs(279) <= not((layer0_outputs(9591)) and (layer0_outputs(3211)));
    layer1_outputs(280) <= not(layer0_outputs(3326));
    layer1_outputs(281) <= not((layer0_outputs(9071)) xor (layer0_outputs(10200)));
    layer1_outputs(282) <= layer0_outputs(9155);
    layer1_outputs(283) <= not((layer0_outputs(3228)) xor (layer0_outputs(3135)));
    layer1_outputs(284) <= not((layer0_outputs(8353)) or (layer0_outputs(1687)));
    layer1_outputs(285) <= layer0_outputs(1119);
    layer1_outputs(286) <= not(layer0_outputs(8282));
    layer1_outputs(287) <= (layer0_outputs(4687)) and not (layer0_outputs(6636));
    layer1_outputs(288) <= not(layer0_outputs(605)) or (layer0_outputs(185));
    layer1_outputs(289) <= (layer0_outputs(4554)) and not (layer0_outputs(4311));
    layer1_outputs(290) <= not(layer0_outputs(9013));
    layer1_outputs(291) <= not(layer0_outputs(5406)) or (layer0_outputs(6977));
    layer1_outputs(292) <= not((layer0_outputs(4860)) or (layer0_outputs(9125)));
    layer1_outputs(293) <= layer0_outputs(10114);
    layer1_outputs(294) <= not((layer0_outputs(7804)) and (layer0_outputs(1068)));
    layer1_outputs(295) <= not(layer0_outputs(2649)) or (layer0_outputs(6027));
    layer1_outputs(296) <= (layer0_outputs(8468)) and not (layer0_outputs(6048));
    layer1_outputs(297) <= layer0_outputs(6900);
    layer1_outputs(298) <= (layer0_outputs(6554)) xor (layer0_outputs(1859));
    layer1_outputs(299) <= layer0_outputs(6933);
    layer1_outputs(300) <= not(layer0_outputs(3202));
    layer1_outputs(301) <= not(layer0_outputs(6321)) or (layer0_outputs(5149));
    layer1_outputs(302) <= (layer0_outputs(8130)) and not (layer0_outputs(6596));
    layer1_outputs(303) <= not((layer0_outputs(4551)) and (layer0_outputs(2974)));
    layer1_outputs(304) <= (layer0_outputs(4819)) and not (layer0_outputs(4449));
    layer1_outputs(305) <= layer0_outputs(4143);
    layer1_outputs(306) <= layer0_outputs(9199);
    layer1_outputs(307) <= not(layer0_outputs(2922));
    layer1_outputs(308) <= not((layer0_outputs(4693)) and (layer0_outputs(645)));
    layer1_outputs(309) <= layer0_outputs(7363);
    layer1_outputs(310) <= not((layer0_outputs(5273)) or (layer0_outputs(4039)));
    layer1_outputs(311) <= (layer0_outputs(5842)) or (layer0_outputs(2328));
    layer1_outputs(312) <= not(layer0_outputs(8152));
    layer1_outputs(313) <= (layer0_outputs(9945)) and not (layer0_outputs(1836));
    layer1_outputs(314) <= not(layer0_outputs(2455));
    layer1_outputs(315) <= (layer0_outputs(3996)) xor (layer0_outputs(7053));
    layer1_outputs(316) <= not(layer0_outputs(1539));
    layer1_outputs(317) <= '1';
    layer1_outputs(318) <= not((layer0_outputs(6699)) or (layer0_outputs(6648)));
    layer1_outputs(319) <= '0';
    layer1_outputs(320) <= not(layer0_outputs(420)) or (layer0_outputs(9087));
    layer1_outputs(321) <= layer0_outputs(3223);
    layer1_outputs(322) <= not(layer0_outputs(9706));
    layer1_outputs(323) <= '0';
    layer1_outputs(324) <= (layer0_outputs(5576)) or (layer0_outputs(6902));
    layer1_outputs(325) <= (layer0_outputs(6477)) or (layer0_outputs(7474));
    layer1_outputs(326) <= (layer0_outputs(8504)) and not (layer0_outputs(7255));
    layer1_outputs(327) <= (layer0_outputs(9688)) and (layer0_outputs(3784));
    layer1_outputs(328) <= not(layer0_outputs(10085));
    layer1_outputs(329) <= '0';
    layer1_outputs(330) <= not((layer0_outputs(3004)) and (layer0_outputs(8996)));
    layer1_outputs(331) <= layer0_outputs(8511);
    layer1_outputs(332) <= (layer0_outputs(3815)) and (layer0_outputs(7529));
    layer1_outputs(333) <= layer0_outputs(4942);
    layer1_outputs(334) <= layer0_outputs(9571);
    layer1_outputs(335) <= (layer0_outputs(7577)) and (layer0_outputs(4291));
    layer1_outputs(336) <= not(layer0_outputs(4007)) or (layer0_outputs(5348));
    layer1_outputs(337) <= layer0_outputs(1613);
    layer1_outputs(338) <= not(layer0_outputs(2662));
    layer1_outputs(339) <= not(layer0_outputs(4643)) or (layer0_outputs(9466));
    layer1_outputs(340) <= not((layer0_outputs(6585)) and (layer0_outputs(357)));
    layer1_outputs(341) <= not(layer0_outputs(126));
    layer1_outputs(342) <= layer0_outputs(8951);
    layer1_outputs(343) <= layer0_outputs(3447);
    layer1_outputs(344) <= layer0_outputs(5107);
    layer1_outputs(345) <= (layer0_outputs(5087)) and not (layer0_outputs(1114));
    layer1_outputs(346) <= (layer0_outputs(7654)) or (layer0_outputs(6460));
    layer1_outputs(347) <= not(layer0_outputs(6087));
    layer1_outputs(348) <= not((layer0_outputs(3593)) and (layer0_outputs(9260)));
    layer1_outputs(349) <= (layer0_outputs(2868)) and not (layer0_outputs(91));
    layer1_outputs(350) <= not(layer0_outputs(2195));
    layer1_outputs(351) <= layer0_outputs(4917);
    layer1_outputs(352) <= '0';
    layer1_outputs(353) <= (layer0_outputs(2383)) or (layer0_outputs(6709));
    layer1_outputs(354) <= not(layer0_outputs(366));
    layer1_outputs(355) <= '0';
    layer1_outputs(356) <= not(layer0_outputs(191));
    layer1_outputs(357) <= '1';
    layer1_outputs(358) <= (layer0_outputs(329)) or (layer0_outputs(9355));
    layer1_outputs(359) <= (layer0_outputs(5380)) and not (layer0_outputs(2632));
    layer1_outputs(360) <= (layer0_outputs(3475)) and not (layer0_outputs(3238));
    layer1_outputs(361) <= (layer0_outputs(1462)) and not (layer0_outputs(7670));
    layer1_outputs(362) <= not(layer0_outputs(9626)) or (layer0_outputs(947));
    layer1_outputs(363) <= '0';
    layer1_outputs(364) <= (layer0_outputs(9878)) xor (layer0_outputs(6087));
    layer1_outputs(365) <= not(layer0_outputs(4246)) or (layer0_outputs(3385));
    layer1_outputs(366) <= not(layer0_outputs(2170));
    layer1_outputs(367) <= (layer0_outputs(1386)) and not (layer0_outputs(6989));
    layer1_outputs(368) <= (layer0_outputs(9802)) or (layer0_outputs(5563));
    layer1_outputs(369) <= not(layer0_outputs(9034)) or (layer0_outputs(3579));
    layer1_outputs(370) <= (layer0_outputs(8089)) and not (layer0_outputs(10039));
    layer1_outputs(371) <= not(layer0_outputs(5048)) or (layer0_outputs(5216));
    layer1_outputs(372) <= (layer0_outputs(2999)) xor (layer0_outputs(6591));
    layer1_outputs(373) <= not(layer0_outputs(6697)) or (layer0_outputs(3540));
    layer1_outputs(374) <= not(layer0_outputs(5311)) or (layer0_outputs(9212));
    layer1_outputs(375) <= not((layer0_outputs(6249)) xor (layer0_outputs(4400)));
    layer1_outputs(376) <= not(layer0_outputs(9352));
    layer1_outputs(377) <= not((layer0_outputs(259)) xor (layer0_outputs(8238)));
    layer1_outputs(378) <= layer0_outputs(9498);
    layer1_outputs(379) <= (layer0_outputs(9443)) and not (layer0_outputs(6931));
    layer1_outputs(380) <= (layer0_outputs(4466)) and not (layer0_outputs(6841));
    layer1_outputs(381) <= not((layer0_outputs(1408)) or (layer0_outputs(4496)));
    layer1_outputs(382) <= not((layer0_outputs(6135)) or (layer0_outputs(1704)));
    layer1_outputs(383) <= (layer0_outputs(7651)) xor (layer0_outputs(7370));
    layer1_outputs(384) <= not((layer0_outputs(8446)) xor (layer0_outputs(1390)));
    layer1_outputs(385) <= not(layer0_outputs(3895));
    layer1_outputs(386) <= (layer0_outputs(606)) and (layer0_outputs(9742));
    layer1_outputs(387) <= layer0_outputs(9294);
    layer1_outputs(388) <= not((layer0_outputs(532)) or (layer0_outputs(6352)));
    layer1_outputs(389) <= not(layer0_outputs(4554));
    layer1_outputs(390) <= layer0_outputs(963);
    layer1_outputs(391) <= layer0_outputs(3706);
    layer1_outputs(392) <= not(layer0_outputs(2006));
    layer1_outputs(393) <= not(layer0_outputs(7131)) or (layer0_outputs(6730));
    layer1_outputs(394) <= layer0_outputs(3059);
    layer1_outputs(395) <= not((layer0_outputs(3513)) or (layer0_outputs(9824)));
    layer1_outputs(396) <= not((layer0_outputs(9366)) xor (layer0_outputs(3013)));
    layer1_outputs(397) <= (layer0_outputs(872)) or (layer0_outputs(771));
    layer1_outputs(398) <= not((layer0_outputs(2544)) and (layer0_outputs(9102)));
    layer1_outputs(399) <= (layer0_outputs(2229)) xor (layer0_outputs(4087));
    layer1_outputs(400) <= not(layer0_outputs(7864)) or (layer0_outputs(4039));
    layer1_outputs(401) <= layer0_outputs(2158);
    layer1_outputs(402) <= layer0_outputs(7790);
    layer1_outputs(403) <= not(layer0_outputs(3855));
    layer1_outputs(404) <= not((layer0_outputs(3024)) xor (layer0_outputs(3780)));
    layer1_outputs(405) <= not(layer0_outputs(3844)) or (layer0_outputs(8380));
    layer1_outputs(406) <= not(layer0_outputs(6017)) or (layer0_outputs(3309));
    layer1_outputs(407) <= (layer0_outputs(3420)) and not (layer0_outputs(4399));
    layer1_outputs(408) <= not(layer0_outputs(3494));
    layer1_outputs(409) <= not((layer0_outputs(779)) and (layer0_outputs(6744)));
    layer1_outputs(410) <= (layer0_outputs(889)) xor (layer0_outputs(4288));
    layer1_outputs(411) <= (layer0_outputs(3748)) and (layer0_outputs(554));
    layer1_outputs(412) <= (layer0_outputs(4990)) and not (layer0_outputs(5931));
    layer1_outputs(413) <= not((layer0_outputs(7382)) xor (layer0_outputs(2130)));
    layer1_outputs(414) <= (layer0_outputs(4989)) xor (layer0_outputs(2740));
    layer1_outputs(415) <= (layer0_outputs(5612)) and not (layer0_outputs(776));
    layer1_outputs(416) <= (layer0_outputs(213)) and not (layer0_outputs(9261));
    layer1_outputs(417) <= not(layer0_outputs(2313));
    layer1_outputs(418) <= (layer0_outputs(7761)) and not (layer0_outputs(7354));
    layer1_outputs(419) <= (layer0_outputs(8584)) and (layer0_outputs(8772));
    layer1_outputs(420) <= (layer0_outputs(8061)) or (layer0_outputs(1775));
    layer1_outputs(421) <= (layer0_outputs(3724)) and not (layer0_outputs(2220));
    layer1_outputs(422) <= not(layer0_outputs(10121)) or (layer0_outputs(1009));
    layer1_outputs(423) <= not((layer0_outputs(5341)) xor (layer0_outputs(1029)));
    layer1_outputs(424) <= layer0_outputs(6128);
    layer1_outputs(425) <= not(layer0_outputs(10035));
    layer1_outputs(426) <= not((layer0_outputs(3084)) or (layer0_outputs(2863)));
    layer1_outputs(427) <= not(layer0_outputs(8317)) or (layer0_outputs(9979));
    layer1_outputs(428) <= not((layer0_outputs(4328)) or (layer0_outputs(8090)));
    layer1_outputs(429) <= layer0_outputs(278);
    layer1_outputs(430) <= layer0_outputs(2354);
    layer1_outputs(431) <= (layer0_outputs(2197)) or (layer0_outputs(4349));
    layer1_outputs(432) <= not(layer0_outputs(233));
    layer1_outputs(433) <= not(layer0_outputs(5897));
    layer1_outputs(434) <= layer0_outputs(2850);
    layer1_outputs(435) <= '0';
    layer1_outputs(436) <= layer0_outputs(782);
    layer1_outputs(437) <= (layer0_outputs(9390)) and (layer0_outputs(2269));
    layer1_outputs(438) <= not((layer0_outputs(4366)) and (layer0_outputs(7022)));
    layer1_outputs(439) <= (layer0_outputs(3201)) and (layer0_outputs(2239));
    layer1_outputs(440) <= (layer0_outputs(2118)) xor (layer0_outputs(4749));
    layer1_outputs(441) <= not((layer0_outputs(3210)) or (layer0_outputs(4572)));
    layer1_outputs(442) <= not(layer0_outputs(160));
    layer1_outputs(443) <= layer0_outputs(8696);
    layer1_outputs(444) <= not((layer0_outputs(2439)) or (layer0_outputs(9278)));
    layer1_outputs(445) <= layer0_outputs(6003);
    layer1_outputs(446) <= not((layer0_outputs(355)) and (layer0_outputs(6425)));
    layer1_outputs(447) <= not(layer0_outputs(7313));
    layer1_outputs(448) <= (layer0_outputs(10081)) xor (layer0_outputs(1599));
    layer1_outputs(449) <= not(layer0_outputs(235));
    layer1_outputs(450) <= not(layer0_outputs(5004)) or (layer0_outputs(8047));
    layer1_outputs(451) <= not(layer0_outputs(6600));
    layer1_outputs(452) <= (layer0_outputs(3936)) and not (layer0_outputs(4732));
    layer1_outputs(453) <= not(layer0_outputs(38));
    layer1_outputs(454) <= not((layer0_outputs(4240)) or (layer0_outputs(757)));
    layer1_outputs(455) <= (layer0_outputs(5183)) and not (layer0_outputs(5459));
    layer1_outputs(456) <= (layer0_outputs(4028)) xor (layer0_outputs(46));
    layer1_outputs(457) <= layer0_outputs(6456);
    layer1_outputs(458) <= not((layer0_outputs(2157)) and (layer0_outputs(4557)));
    layer1_outputs(459) <= layer0_outputs(116);
    layer1_outputs(460) <= (layer0_outputs(2050)) and not (layer0_outputs(9151));
    layer1_outputs(461) <= not((layer0_outputs(6180)) or (layer0_outputs(3505)));
    layer1_outputs(462) <= layer0_outputs(9350);
    layer1_outputs(463) <= not(layer0_outputs(4787)) or (layer0_outputs(7730));
    layer1_outputs(464) <= (layer0_outputs(3952)) and (layer0_outputs(6507));
    layer1_outputs(465) <= not(layer0_outputs(9699)) or (layer0_outputs(3825));
    layer1_outputs(466) <= not(layer0_outputs(8162));
    layer1_outputs(467) <= not((layer0_outputs(7312)) and (layer0_outputs(3775)));
    layer1_outputs(468) <= (layer0_outputs(7928)) and (layer0_outputs(6380));
    layer1_outputs(469) <= not(layer0_outputs(2167)) or (layer0_outputs(9908));
    layer1_outputs(470) <= (layer0_outputs(3764)) and (layer0_outputs(4943));
    layer1_outputs(471) <= (layer0_outputs(7466)) or (layer0_outputs(10024));
    layer1_outputs(472) <= layer0_outputs(5658);
    layer1_outputs(473) <= layer0_outputs(2343);
    layer1_outputs(474) <= layer0_outputs(9202);
    layer1_outputs(475) <= not(layer0_outputs(8794)) or (layer0_outputs(7605));
    layer1_outputs(476) <= (layer0_outputs(7007)) and not (layer0_outputs(8471));
    layer1_outputs(477) <= not(layer0_outputs(9036));
    layer1_outputs(478) <= (layer0_outputs(6227)) xor (layer0_outputs(3954));
    layer1_outputs(479) <= not((layer0_outputs(9196)) and (layer0_outputs(398)));
    layer1_outputs(480) <= (layer0_outputs(1773)) and not (layer0_outputs(6654));
    layer1_outputs(481) <= (layer0_outputs(4684)) xor (layer0_outputs(7696));
    layer1_outputs(482) <= (layer0_outputs(7759)) or (layer0_outputs(4782));
    layer1_outputs(483) <= not(layer0_outputs(279));
    layer1_outputs(484) <= (layer0_outputs(3482)) and not (layer0_outputs(4736));
    layer1_outputs(485) <= not(layer0_outputs(2130)) or (layer0_outputs(3269));
    layer1_outputs(486) <= not(layer0_outputs(4856));
    layer1_outputs(487) <= (layer0_outputs(1645)) xor (layer0_outputs(6686));
    layer1_outputs(488) <= not((layer0_outputs(6852)) and (layer0_outputs(8196)));
    layer1_outputs(489) <= not(layer0_outputs(2129));
    layer1_outputs(490) <= not(layer0_outputs(7935)) or (layer0_outputs(9717));
    layer1_outputs(491) <= (layer0_outputs(2067)) and not (layer0_outputs(5088));
    layer1_outputs(492) <= not(layer0_outputs(2925)) or (layer0_outputs(1138));
    layer1_outputs(493) <= (layer0_outputs(7960)) and (layer0_outputs(4717));
    layer1_outputs(494) <= not(layer0_outputs(2676));
    layer1_outputs(495) <= layer0_outputs(8007);
    layer1_outputs(496) <= (layer0_outputs(1132)) and not (layer0_outputs(7025));
    layer1_outputs(497) <= not(layer0_outputs(3139));
    layer1_outputs(498) <= not(layer0_outputs(868)) or (layer0_outputs(761));
    layer1_outputs(499) <= '0';
    layer1_outputs(500) <= layer0_outputs(4328);
    layer1_outputs(501) <= not((layer0_outputs(174)) and (layer0_outputs(5291)));
    layer1_outputs(502) <= (layer0_outputs(2609)) and (layer0_outputs(6671));
    layer1_outputs(503) <= layer0_outputs(2006);
    layer1_outputs(504) <= not(layer0_outputs(10059));
    layer1_outputs(505) <= layer0_outputs(5639);
    layer1_outputs(506) <= layer0_outputs(5393);
    layer1_outputs(507) <= not(layer0_outputs(3427)) or (layer0_outputs(9117));
    layer1_outputs(508) <= not((layer0_outputs(5209)) and (layer0_outputs(5854)));
    layer1_outputs(509) <= (layer0_outputs(4536)) xor (layer0_outputs(5285));
    layer1_outputs(510) <= (layer0_outputs(8104)) and not (layer0_outputs(825));
    layer1_outputs(511) <= (layer0_outputs(6915)) and not (layer0_outputs(1594));
    layer1_outputs(512) <= (layer0_outputs(529)) and (layer0_outputs(10048));
    layer1_outputs(513) <= (layer0_outputs(2346)) xor (layer0_outputs(8214));
    layer1_outputs(514) <= (layer0_outputs(5399)) xor (layer0_outputs(7337));
    layer1_outputs(515) <= layer0_outputs(3555);
    layer1_outputs(516) <= not((layer0_outputs(6894)) xor (layer0_outputs(9860)));
    layer1_outputs(517) <= (layer0_outputs(7344)) and not (layer0_outputs(1888));
    layer1_outputs(518) <= not(layer0_outputs(8671)) or (layer0_outputs(4258));
    layer1_outputs(519) <= layer0_outputs(8475);
    layer1_outputs(520) <= not(layer0_outputs(5841)) or (layer0_outputs(6950));
    layer1_outputs(521) <= layer0_outputs(1324);
    layer1_outputs(522) <= not(layer0_outputs(4478));
    layer1_outputs(523) <= not(layer0_outputs(7830)) or (layer0_outputs(15));
    layer1_outputs(524) <= (layer0_outputs(2104)) and (layer0_outputs(6027));
    layer1_outputs(525) <= (layer0_outputs(7543)) and (layer0_outputs(7856));
    layer1_outputs(526) <= (layer0_outputs(1065)) and not (layer0_outputs(8638));
    layer1_outputs(527) <= not(layer0_outputs(3115));
    layer1_outputs(528) <= not((layer0_outputs(8912)) or (layer0_outputs(2441)));
    layer1_outputs(529) <= not((layer0_outputs(9181)) xor (layer0_outputs(8947)));
    layer1_outputs(530) <= (layer0_outputs(5779)) xor (layer0_outputs(8674));
    layer1_outputs(531) <= (layer0_outputs(2180)) and not (layer0_outputs(7579));
    layer1_outputs(532) <= not((layer0_outputs(8244)) xor (layer0_outputs(5047)));
    layer1_outputs(533) <= not(layer0_outputs(5986)) or (layer0_outputs(3658));
    layer1_outputs(534) <= not((layer0_outputs(5489)) or (layer0_outputs(4295)));
    layer1_outputs(535) <= (layer0_outputs(5174)) xor (layer0_outputs(2136));
    layer1_outputs(536) <= not(layer0_outputs(5463));
    layer1_outputs(537) <= not(layer0_outputs(5172));
    layer1_outputs(538) <= layer0_outputs(2588);
    layer1_outputs(539) <= layer0_outputs(7325);
    layer1_outputs(540) <= not(layer0_outputs(5592));
    layer1_outputs(541) <= '1';
    layer1_outputs(542) <= layer0_outputs(6300);
    layer1_outputs(543) <= '0';
    layer1_outputs(544) <= not(layer0_outputs(7402)) or (layer0_outputs(5254));
    layer1_outputs(545) <= layer0_outputs(2584);
    layer1_outputs(546) <= not((layer0_outputs(6707)) or (layer0_outputs(7712)));
    layer1_outputs(547) <= not(layer0_outputs(10064));
    layer1_outputs(548) <= (layer0_outputs(5916)) or (layer0_outputs(7793));
    layer1_outputs(549) <= layer0_outputs(8406);
    layer1_outputs(550) <= not(layer0_outputs(2603));
    layer1_outputs(551) <= layer0_outputs(539);
    layer1_outputs(552) <= not(layer0_outputs(9363));
    layer1_outputs(553) <= (layer0_outputs(7273)) or (layer0_outputs(8974));
    layer1_outputs(554) <= (layer0_outputs(2895)) xor (layer0_outputs(8163));
    layer1_outputs(555) <= (layer0_outputs(8719)) xor (layer0_outputs(19));
    layer1_outputs(556) <= not((layer0_outputs(5096)) or (layer0_outputs(1059)));
    layer1_outputs(557) <= not(layer0_outputs(273)) or (layer0_outputs(6838));
    layer1_outputs(558) <= not((layer0_outputs(3524)) or (layer0_outputs(4708)));
    layer1_outputs(559) <= (layer0_outputs(7844)) xor (layer0_outputs(4747));
    layer1_outputs(560) <= (layer0_outputs(5891)) and not (layer0_outputs(6517));
    layer1_outputs(561) <= not(layer0_outputs(8982)) or (layer0_outputs(9379));
    layer1_outputs(562) <= not(layer0_outputs(5238));
    layer1_outputs(563) <= layer0_outputs(4063);
    layer1_outputs(564) <= (layer0_outputs(9691)) and not (layer0_outputs(544));
    layer1_outputs(565) <= (layer0_outputs(9032)) and not (layer0_outputs(5579));
    layer1_outputs(566) <= layer0_outputs(2375);
    layer1_outputs(567) <= not((layer0_outputs(5583)) xor (layer0_outputs(6071)));
    layer1_outputs(568) <= not(layer0_outputs(7536));
    layer1_outputs(569) <= not((layer0_outputs(1942)) xor (layer0_outputs(9559)));
    layer1_outputs(570) <= '1';
    layer1_outputs(571) <= not(layer0_outputs(7166));
    layer1_outputs(572) <= (layer0_outputs(6823)) xor (layer0_outputs(2878));
    layer1_outputs(573) <= (layer0_outputs(6888)) or (layer0_outputs(9103));
    layer1_outputs(574) <= (layer0_outputs(8091)) and (layer0_outputs(7490));
    layer1_outputs(575) <= not(layer0_outputs(1864));
    layer1_outputs(576) <= not(layer0_outputs(1907));
    layer1_outputs(577) <= not(layer0_outputs(3059));
    layer1_outputs(578) <= not(layer0_outputs(6514)) or (layer0_outputs(6628));
    layer1_outputs(579) <= layer0_outputs(8275);
    layer1_outputs(580) <= layer0_outputs(7770);
    layer1_outputs(581) <= not(layer0_outputs(3793));
    layer1_outputs(582) <= not(layer0_outputs(8234)) or (layer0_outputs(2386));
    layer1_outputs(583) <= layer0_outputs(6786);
    layer1_outputs(584) <= not((layer0_outputs(4920)) or (layer0_outputs(2971)));
    layer1_outputs(585) <= layer0_outputs(4994);
    layer1_outputs(586) <= layer0_outputs(7734);
    layer1_outputs(587) <= layer0_outputs(9518);
    layer1_outputs(588) <= (layer0_outputs(269)) and not (layer0_outputs(5180));
    layer1_outputs(589) <= (layer0_outputs(6807)) and (layer0_outputs(283));
    layer1_outputs(590) <= (layer0_outputs(6564)) and not (layer0_outputs(4031));
    layer1_outputs(591) <= (layer0_outputs(1792)) xor (layer0_outputs(3632));
    layer1_outputs(592) <= layer0_outputs(6186);
    layer1_outputs(593) <= not(layer0_outputs(1680)) or (layer0_outputs(4278));
    layer1_outputs(594) <= not((layer0_outputs(6199)) or (layer0_outputs(8395)));
    layer1_outputs(595) <= not(layer0_outputs(5966));
    layer1_outputs(596) <= (layer0_outputs(9369)) or (layer0_outputs(2950));
    layer1_outputs(597) <= (layer0_outputs(3209)) or (layer0_outputs(9757));
    layer1_outputs(598) <= not((layer0_outputs(8753)) or (layer0_outputs(2377)));
    layer1_outputs(599) <= '1';
    layer1_outputs(600) <= not(layer0_outputs(6395));
    layer1_outputs(601) <= (layer0_outputs(7134)) xor (layer0_outputs(368));
    layer1_outputs(602) <= (layer0_outputs(4204)) and (layer0_outputs(9100));
    layer1_outputs(603) <= not(layer0_outputs(3245)) or (layer0_outputs(4223));
    layer1_outputs(604) <= (layer0_outputs(9810)) xor (layer0_outputs(9697));
    layer1_outputs(605) <= (layer0_outputs(8673)) or (layer0_outputs(10075));
    layer1_outputs(606) <= layer0_outputs(3074);
    layer1_outputs(607) <= (layer0_outputs(5724)) or (layer0_outputs(7088));
    layer1_outputs(608) <= not(layer0_outputs(5106)) or (layer0_outputs(5635));
    layer1_outputs(609) <= (layer0_outputs(3240)) and not (layer0_outputs(7454));
    layer1_outputs(610) <= not(layer0_outputs(711));
    layer1_outputs(611) <= not((layer0_outputs(9420)) xor (layer0_outputs(10092)));
    layer1_outputs(612) <= not((layer0_outputs(5959)) xor (layer0_outputs(4974)));
    layer1_outputs(613) <= not(layer0_outputs(688)) or (layer0_outputs(828));
    layer1_outputs(614) <= layer0_outputs(391);
    layer1_outputs(615) <= (layer0_outputs(4627)) and not (layer0_outputs(4133));
    layer1_outputs(616) <= not(layer0_outputs(7381));
    layer1_outputs(617) <= layer0_outputs(3535);
    layer1_outputs(618) <= layer0_outputs(9316);
    layer1_outputs(619) <= layer0_outputs(1408);
    layer1_outputs(620) <= (layer0_outputs(7200)) or (layer0_outputs(1116));
    layer1_outputs(621) <= not(layer0_outputs(3323)) or (layer0_outputs(7647));
    layer1_outputs(622) <= not(layer0_outputs(9335)) or (layer0_outputs(9481));
    layer1_outputs(623) <= not(layer0_outputs(4893));
    layer1_outputs(624) <= (layer0_outputs(281)) and (layer0_outputs(721));
    layer1_outputs(625) <= (layer0_outputs(5603)) and not (layer0_outputs(1947));
    layer1_outputs(626) <= not(layer0_outputs(4236));
    layer1_outputs(627) <= not((layer0_outputs(7590)) xor (layer0_outputs(7823)));
    layer1_outputs(628) <= not(layer0_outputs(110));
    layer1_outputs(629) <= not(layer0_outputs(4739));
    layer1_outputs(630) <= (layer0_outputs(7987)) and not (layer0_outputs(8847));
    layer1_outputs(631) <= layer0_outputs(1790);
    layer1_outputs(632) <= layer0_outputs(8718);
    layer1_outputs(633) <= layer0_outputs(10171);
    layer1_outputs(634) <= not(layer0_outputs(7495));
    layer1_outputs(635) <= not((layer0_outputs(1620)) and (layer0_outputs(514)));
    layer1_outputs(636) <= not(layer0_outputs(2094)) or (layer0_outputs(5551));
    layer1_outputs(637) <= (layer0_outputs(2637)) or (layer0_outputs(4999));
    layer1_outputs(638) <= (layer0_outputs(7414)) xor (layer0_outputs(604));
    layer1_outputs(639) <= not((layer0_outputs(7888)) and (layer0_outputs(744)));
    layer1_outputs(640) <= layer0_outputs(7709);
    layer1_outputs(641) <= '1';
    layer1_outputs(642) <= layer0_outputs(4512);
    layer1_outputs(643) <= layer0_outputs(1195);
    layer1_outputs(644) <= not(layer0_outputs(536));
    layer1_outputs(645) <= not((layer0_outputs(80)) xor (layer0_outputs(9448)));
    layer1_outputs(646) <= not(layer0_outputs(7058));
    layer1_outputs(647) <= not((layer0_outputs(7050)) or (layer0_outputs(9104)));
    layer1_outputs(648) <= not(layer0_outputs(3302));
    layer1_outputs(649) <= (layer0_outputs(5511)) or (layer0_outputs(3206));
    layer1_outputs(650) <= not(layer0_outputs(2355));
    layer1_outputs(651) <= (layer0_outputs(7410)) and (layer0_outputs(8566));
    layer1_outputs(652) <= not(layer0_outputs(2743));
    layer1_outputs(653) <= (layer0_outputs(9651)) or (layer0_outputs(7578));
    layer1_outputs(654) <= not((layer0_outputs(9451)) or (layer0_outputs(8236)));
    layer1_outputs(655) <= (layer0_outputs(6915)) and (layer0_outputs(785));
    layer1_outputs(656) <= not(layer0_outputs(6677));
    layer1_outputs(657) <= (layer0_outputs(7621)) and (layer0_outputs(7491));
    layer1_outputs(658) <= not(layer0_outputs(5913));
    layer1_outputs(659) <= layer0_outputs(369);
    layer1_outputs(660) <= layer0_outputs(9123);
    layer1_outputs(661) <= (layer0_outputs(331)) xor (layer0_outputs(5148));
    layer1_outputs(662) <= layer0_outputs(1997);
    layer1_outputs(663) <= layer0_outputs(8797);
    layer1_outputs(664) <= not(layer0_outputs(1603)) or (layer0_outputs(3382));
    layer1_outputs(665) <= (layer0_outputs(4256)) xor (layer0_outputs(8335));
    layer1_outputs(666) <= (layer0_outputs(5123)) and (layer0_outputs(6063));
    layer1_outputs(667) <= not((layer0_outputs(6300)) and (layer0_outputs(5866)));
    layer1_outputs(668) <= not(layer0_outputs(3972)) or (layer0_outputs(4520));
    layer1_outputs(669) <= (layer0_outputs(6986)) and (layer0_outputs(706));
    layer1_outputs(670) <= (layer0_outputs(2143)) and not (layer0_outputs(2810));
    layer1_outputs(671) <= layer0_outputs(4189);
    layer1_outputs(672) <= (layer0_outputs(2029)) and not (layer0_outputs(5108));
    layer1_outputs(673) <= (layer0_outputs(7491)) and not (layer0_outputs(8789));
    layer1_outputs(674) <= not((layer0_outputs(9028)) xor (layer0_outputs(7779)));
    layer1_outputs(675) <= (layer0_outputs(953)) and (layer0_outputs(4591));
    layer1_outputs(676) <= (layer0_outputs(3343)) and not (layer0_outputs(7195));
    layer1_outputs(677) <= not(layer0_outputs(6207));
    layer1_outputs(678) <= not(layer0_outputs(8725)) or (layer0_outputs(8357));
    layer1_outputs(679) <= (layer0_outputs(7597)) or (layer0_outputs(9053));
    layer1_outputs(680) <= layer0_outputs(4055);
    layer1_outputs(681) <= not(layer0_outputs(5471));
    layer1_outputs(682) <= (layer0_outputs(1345)) xor (layer0_outputs(1520));
    layer1_outputs(683) <= not(layer0_outputs(2511));
    layer1_outputs(684) <= not(layer0_outputs(1139));
    layer1_outputs(685) <= not(layer0_outputs(5178));
    layer1_outputs(686) <= not(layer0_outputs(9973)) or (layer0_outputs(7240));
    layer1_outputs(687) <= not(layer0_outputs(39));
    layer1_outputs(688) <= layer0_outputs(2012);
    layer1_outputs(689) <= not(layer0_outputs(1755));
    layer1_outputs(690) <= not(layer0_outputs(9128));
    layer1_outputs(691) <= not(layer0_outputs(1611));
    layer1_outputs(692) <= layer0_outputs(665);
    layer1_outputs(693) <= layer0_outputs(6917);
    layer1_outputs(694) <= '1';
    layer1_outputs(695) <= (layer0_outputs(2139)) and not (layer0_outputs(9412));
    layer1_outputs(696) <= (layer0_outputs(3029)) or (layer0_outputs(8175));
    layer1_outputs(697) <= layer0_outputs(1206);
    layer1_outputs(698) <= (layer0_outputs(2192)) and not (layer0_outputs(1828));
    layer1_outputs(699) <= (layer0_outputs(1612)) and (layer0_outputs(1251));
    layer1_outputs(700) <= not(layer0_outputs(1064)) or (layer0_outputs(7867));
    layer1_outputs(701) <= not((layer0_outputs(2794)) or (layer0_outputs(2972)));
    layer1_outputs(702) <= layer0_outputs(8321);
    layer1_outputs(703) <= (layer0_outputs(6257)) and (layer0_outputs(479));
    layer1_outputs(704) <= not(layer0_outputs(2350));
    layer1_outputs(705) <= not((layer0_outputs(4845)) or (layer0_outputs(4552)));
    layer1_outputs(706) <= not(layer0_outputs(3584)) or (layer0_outputs(3085));
    layer1_outputs(707) <= not((layer0_outputs(1405)) or (layer0_outputs(8027)));
    layer1_outputs(708) <= not(layer0_outputs(6007)) or (layer0_outputs(627));
    layer1_outputs(709) <= (layer0_outputs(988)) and not (layer0_outputs(183));
    layer1_outputs(710) <= not((layer0_outputs(3495)) and (layer0_outputs(4231)));
    layer1_outputs(711) <= not(layer0_outputs(1483));
    layer1_outputs(712) <= not(layer0_outputs(6684));
    layer1_outputs(713) <= not((layer0_outputs(2311)) and (layer0_outputs(6305)));
    layer1_outputs(714) <= not(layer0_outputs(4575));
    layer1_outputs(715) <= (layer0_outputs(1058)) and (layer0_outputs(1860));
    layer1_outputs(716) <= not(layer0_outputs(1551)) or (layer0_outputs(2359));
    layer1_outputs(717) <= '0';
    layer1_outputs(718) <= (layer0_outputs(10167)) xor (layer0_outputs(9469));
    layer1_outputs(719) <= not((layer0_outputs(7359)) or (layer0_outputs(2850)));
    layer1_outputs(720) <= '1';
    layer1_outputs(721) <= layer0_outputs(3514);
    layer1_outputs(722) <= layer0_outputs(7632);
    layer1_outputs(723) <= not(layer0_outputs(2309));
    layer1_outputs(724) <= not(layer0_outputs(2068));
    layer1_outputs(725) <= not((layer0_outputs(2519)) or (layer0_outputs(3674)));
    layer1_outputs(726) <= not((layer0_outputs(6445)) and (layer0_outputs(8837)));
    layer1_outputs(727) <= not(layer0_outputs(5954)) or (layer0_outputs(8426));
    layer1_outputs(728) <= layer0_outputs(8628);
    layer1_outputs(729) <= (layer0_outputs(7985)) and (layer0_outputs(1371));
    layer1_outputs(730) <= layer0_outputs(2152);
    layer1_outputs(731) <= (layer0_outputs(1053)) and not (layer0_outputs(3796));
    layer1_outputs(732) <= not((layer0_outputs(2663)) xor (layer0_outputs(1764)));
    layer1_outputs(733) <= not(layer0_outputs(2288));
    layer1_outputs(734) <= (layer0_outputs(4765)) and not (layer0_outputs(8836));
    layer1_outputs(735) <= (layer0_outputs(694)) and (layer0_outputs(9819));
    layer1_outputs(736) <= '0';
    layer1_outputs(737) <= (layer0_outputs(3877)) and not (layer0_outputs(4965));
    layer1_outputs(738) <= not((layer0_outputs(3978)) and (layer0_outputs(3159)));
    layer1_outputs(739) <= (layer0_outputs(8903)) or (layer0_outputs(2662));
    layer1_outputs(740) <= not(layer0_outputs(75)) or (layer0_outputs(9701));
    layer1_outputs(741) <= not((layer0_outputs(298)) and (layer0_outputs(10009)));
    layer1_outputs(742) <= (layer0_outputs(5250)) xor (layer0_outputs(2186));
    layer1_outputs(743) <= '1';
    layer1_outputs(744) <= not((layer0_outputs(1235)) or (layer0_outputs(892)));
    layer1_outputs(745) <= layer0_outputs(2182);
    layer1_outputs(746) <= layer0_outputs(4216);
    layer1_outputs(747) <= '0';
    layer1_outputs(748) <= (layer0_outputs(1380)) and not (layer0_outputs(8679));
    layer1_outputs(749) <= not((layer0_outputs(2875)) xor (layer0_outputs(1331)));
    layer1_outputs(750) <= not(layer0_outputs(8203));
    layer1_outputs(751) <= (layer0_outputs(373)) and not (layer0_outputs(7366));
    layer1_outputs(752) <= (layer0_outputs(3615)) or (layer0_outputs(360));
    layer1_outputs(753) <= not((layer0_outputs(6)) xor (layer0_outputs(8989)));
    layer1_outputs(754) <= (layer0_outputs(21)) and not (layer0_outputs(6047));
    layer1_outputs(755) <= not(layer0_outputs(4272));
    layer1_outputs(756) <= (layer0_outputs(10090)) and (layer0_outputs(5616));
    layer1_outputs(757) <= (layer0_outputs(948)) and not (layer0_outputs(8031));
    layer1_outputs(758) <= (layer0_outputs(8795)) or (layer0_outputs(6090));
    layer1_outputs(759) <= not(layer0_outputs(8968));
    layer1_outputs(760) <= not((layer0_outputs(6330)) or (layer0_outputs(4219)));
    layer1_outputs(761) <= layer0_outputs(5418);
    layer1_outputs(762) <= (layer0_outputs(1623)) and not (layer0_outputs(552));
    layer1_outputs(763) <= (layer0_outputs(7203)) and not (layer0_outputs(57));
    layer1_outputs(764) <= (layer0_outputs(8255)) xor (layer0_outputs(8586));
    layer1_outputs(765) <= not(layer0_outputs(1654));
    layer1_outputs(766) <= (layer0_outputs(3010)) and not (layer0_outputs(7948));
    layer1_outputs(767) <= not(layer0_outputs(3346)) or (layer0_outputs(8804));
    layer1_outputs(768) <= not(layer0_outputs(1017));
    layer1_outputs(769) <= not(layer0_outputs(8719));
    layer1_outputs(770) <= (layer0_outputs(3170)) or (layer0_outputs(7879));
    layer1_outputs(771) <= layer0_outputs(9484);
    layer1_outputs(772) <= not(layer0_outputs(3839)) or (layer0_outputs(7993));
    layer1_outputs(773) <= layer0_outputs(3860);
    layer1_outputs(774) <= not(layer0_outputs(6889));
    layer1_outputs(775) <= not(layer0_outputs(1043));
    layer1_outputs(776) <= layer0_outputs(1574);
    layer1_outputs(777) <= layer0_outputs(3414);
    layer1_outputs(778) <= layer0_outputs(5862);
    layer1_outputs(779) <= layer0_outputs(2127);
    layer1_outputs(780) <= (layer0_outputs(3364)) xor (layer0_outputs(1209));
    layer1_outputs(781) <= '0';
    layer1_outputs(782) <= layer0_outputs(5601);
    layer1_outputs(783) <= not(layer0_outputs(214)) or (layer0_outputs(5222));
    layer1_outputs(784) <= not(layer0_outputs(4404));
    layer1_outputs(785) <= (layer0_outputs(6011)) or (layer0_outputs(4410));
    layer1_outputs(786) <= (layer0_outputs(197)) or (layer0_outputs(1365));
    layer1_outputs(787) <= (layer0_outputs(5027)) or (layer0_outputs(6356));
    layer1_outputs(788) <= not(layer0_outputs(5037));
    layer1_outputs(789) <= layer0_outputs(3226);
    layer1_outputs(790) <= layer0_outputs(7925);
    layer1_outputs(791) <= layer0_outputs(7693);
    layer1_outputs(792) <= not(layer0_outputs(7460));
    layer1_outputs(793) <= layer0_outputs(327);
    layer1_outputs(794) <= not((layer0_outputs(4183)) or (layer0_outputs(8022)));
    layer1_outputs(795) <= layer0_outputs(6801);
    layer1_outputs(796) <= not(layer0_outputs(6961));
    layer1_outputs(797) <= not(layer0_outputs(3182)) or (layer0_outputs(591));
    layer1_outputs(798) <= not(layer0_outputs(7214)) or (layer0_outputs(9116));
    layer1_outputs(799) <= layer0_outputs(1878);
    layer1_outputs(800) <= (layer0_outputs(565)) or (layer0_outputs(1616));
    layer1_outputs(801) <= not(layer0_outputs(1363)) or (layer0_outputs(3636));
    layer1_outputs(802) <= layer0_outputs(9960);
    layer1_outputs(803) <= (layer0_outputs(380)) and (layer0_outputs(4834));
    layer1_outputs(804) <= not(layer0_outputs(2368)) or (layer0_outputs(5345));
    layer1_outputs(805) <= layer0_outputs(8712);
    layer1_outputs(806) <= not(layer0_outputs(5653));
    layer1_outputs(807) <= (layer0_outputs(3243)) and not (layer0_outputs(1222));
    layer1_outputs(808) <= layer0_outputs(3906);
    layer1_outputs(809) <= not(layer0_outputs(8383));
    layer1_outputs(810) <= (layer0_outputs(6188)) or (layer0_outputs(2586));
    layer1_outputs(811) <= layer0_outputs(1581);
    layer1_outputs(812) <= layer0_outputs(4549);
    layer1_outputs(813) <= (layer0_outputs(801)) and (layer0_outputs(2802));
    layer1_outputs(814) <= not(layer0_outputs(6213));
    layer1_outputs(815) <= (layer0_outputs(7092)) and (layer0_outputs(4158));
    layer1_outputs(816) <= (layer0_outputs(1051)) and not (layer0_outputs(274));
    layer1_outputs(817) <= not(layer0_outputs(9584));
    layer1_outputs(818) <= (layer0_outputs(2570)) xor (layer0_outputs(9688));
    layer1_outputs(819) <= layer0_outputs(4811);
    layer1_outputs(820) <= not(layer0_outputs(5355));
    layer1_outputs(821) <= (layer0_outputs(7123)) or (layer0_outputs(1925));
    layer1_outputs(822) <= not((layer0_outputs(1763)) xor (layer0_outputs(8579)));
    layer1_outputs(823) <= layer0_outputs(1343);
    layer1_outputs(824) <= layer0_outputs(9239);
    layer1_outputs(825) <= (layer0_outputs(9424)) and not (layer0_outputs(5626));
    layer1_outputs(826) <= (layer0_outputs(4665)) xor (layer0_outputs(3914));
    layer1_outputs(827) <= (layer0_outputs(2834)) or (layer0_outputs(1239));
    layer1_outputs(828) <= layer0_outputs(4899);
    layer1_outputs(829) <= layer0_outputs(156);
    layer1_outputs(830) <= '0';
    layer1_outputs(831) <= (layer0_outputs(7027)) and not (layer0_outputs(4574));
    layer1_outputs(832) <= not(layer0_outputs(9002));
    layer1_outputs(833) <= (layer0_outputs(3560)) and not (layer0_outputs(3645));
    layer1_outputs(834) <= (layer0_outputs(1133)) xor (layer0_outputs(200));
    layer1_outputs(835) <= layer0_outputs(5123);
    layer1_outputs(836) <= (layer0_outputs(6037)) and not (layer0_outputs(3880));
    layer1_outputs(837) <= '1';
    layer1_outputs(838) <= layer0_outputs(4072);
    layer1_outputs(839) <= (layer0_outputs(6811)) and not (layer0_outputs(2550));
    layer1_outputs(840) <= not(layer0_outputs(5366)) or (layer0_outputs(6975));
    layer1_outputs(841) <= layer0_outputs(2171);
    layer1_outputs(842) <= (layer0_outputs(9058)) xor (layer0_outputs(9662));
    layer1_outputs(843) <= not((layer0_outputs(1145)) and (layer0_outputs(6728)));
    layer1_outputs(844) <= not((layer0_outputs(8174)) xor (layer0_outputs(7941)));
    layer1_outputs(845) <= layer0_outputs(6112);
    layer1_outputs(846) <= not(layer0_outputs(655));
    layer1_outputs(847) <= (layer0_outputs(9560)) and (layer0_outputs(4632));
    layer1_outputs(848) <= not(layer0_outputs(4469)) or (layer0_outputs(9216));
    layer1_outputs(849) <= layer0_outputs(7841);
    layer1_outputs(850) <= (layer0_outputs(9936)) and not (layer0_outputs(8360));
    layer1_outputs(851) <= not(layer0_outputs(7726));
    layer1_outputs(852) <= layer0_outputs(5340);
    layer1_outputs(853) <= (layer0_outputs(9580)) and (layer0_outputs(5456));
    layer1_outputs(854) <= not(layer0_outputs(5081));
    layer1_outputs(855) <= not(layer0_outputs(7427)) or (layer0_outputs(2257));
    layer1_outputs(856) <= (layer0_outputs(6527)) and not (layer0_outputs(6264));
    layer1_outputs(857) <= (layer0_outputs(6085)) and not (layer0_outputs(9171));
    layer1_outputs(858) <= (layer0_outputs(4102)) xor (layer0_outputs(7484));
    layer1_outputs(859) <= layer0_outputs(7429);
    layer1_outputs(860) <= (layer0_outputs(2302)) xor (layer0_outputs(5978));
    layer1_outputs(861) <= layer0_outputs(5282);
    layer1_outputs(862) <= not((layer0_outputs(2044)) xor (layer0_outputs(7084)));
    layer1_outputs(863) <= not((layer0_outputs(9634)) and (layer0_outputs(9867)));
    layer1_outputs(864) <= not((layer0_outputs(6113)) and (layer0_outputs(3653)));
    layer1_outputs(865) <= not(layer0_outputs(6803));
    layer1_outputs(866) <= not((layer0_outputs(555)) and (layer0_outputs(8862)));
    layer1_outputs(867) <= not(layer0_outputs(5235));
    layer1_outputs(868) <= not((layer0_outputs(2753)) and (layer0_outputs(9015)));
    layer1_outputs(869) <= (layer0_outputs(1639)) or (layer0_outputs(289));
    layer1_outputs(870) <= not(layer0_outputs(7496));
    layer1_outputs(871) <= not((layer0_outputs(8325)) or (layer0_outputs(8108)));
    layer1_outputs(872) <= '1';
    layer1_outputs(873) <= (layer0_outputs(466)) and not (layer0_outputs(5297));
    layer1_outputs(874) <= not(layer0_outputs(2075));
    layer1_outputs(875) <= not((layer0_outputs(6083)) and (layer0_outputs(5842)));
    layer1_outputs(876) <= not(layer0_outputs(6442));
    layer1_outputs(877) <= not(layer0_outputs(5395)) or (layer0_outputs(9109));
    layer1_outputs(878) <= not((layer0_outputs(1752)) or (layer0_outputs(9349)));
    layer1_outputs(879) <= not(layer0_outputs(1820));
    layer1_outputs(880) <= (layer0_outputs(3448)) and (layer0_outputs(1019));
    layer1_outputs(881) <= not(layer0_outputs(9951));
    layer1_outputs(882) <= (layer0_outputs(1033)) and (layer0_outputs(9988));
    layer1_outputs(883) <= (layer0_outputs(9725)) and not (layer0_outputs(4864));
    layer1_outputs(884) <= not((layer0_outputs(8611)) and (layer0_outputs(3619)));
    layer1_outputs(885) <= not(layer0_outputs(844));
    layer1_outputs(886) <= not(layer0_outputs(3087)) or (layer0_outputs(3695));
    layer1_outputs(887) <= not(layer0_outputs(1227)) or (layer0_outputs(2518));
    layer1_outputs(888) <= (layer0_outputs(2826)) or (layer0_outputs(1491));
    layer1_outputs(889) <= not((layer0_outputs(6883)) xor (layer0_outputs(1248)));
    layer1_outputs(890) <= (layer0_outputs(1881)) or (layer0_outputs(10103));
    layer1_outputs(891) <= not(layer0_outputs(3937));
    layer1_outputs(892) <= (layer0_outputs(5327)) and not (layer0_outputs(9995));
    layer1_outputs(893) <= layer0_outputs(3955);
    layer1_outputs(894) <= not(layer0_outputs(8560));
    layer1_outputs(895) <= (layer0_outputs(1205)) or (layer0_outputs(8698));
    layer1_outputs(896) <= layer0_outputs(9568);
    layer1_outputs(897) <= not(layer0_outputs(5639)) or (layer0_outputs(500));
    layer1_outputs(898) <= layer0_outputs(9568);
    layer1_outputs(899) <= not(layer0_outputs(7552)) or (layer0_outputs(9150));
    layer1_outputs(900) <= not(layer0_outputs(1816)) or (layer0_outputs(2485));
    layer1_outputs(901) <= (layer0_outputs(7371)) and not (layer0_outputs(1858));
    layer1_outputs(902) <= not(layer0_outputs(3137));
    layer1_outputs(903) <= (layer0_outputs(3609)) and not (layer0_outputs(8481));
    layer1_outputs(904) <= '0';
    layer1_outputs(905) <= not(layer0_outputs(240)) or (layer0_outputs(4242));
    layer1_outputs(906) <= layer0_outputs(7589);
    layer1_outputs(907) <= (layer0_outputs(8005)) or (layer0_outputs(6498));
    layer1_outputs(908) <= not(layer0_outputs(4045)) or (layer0_outputs(7202));
    layer1_outputs(909) <= (layer0_outputs(8640)) and (layer0_outputs(7991));
    layer1_outputs(910) <= not(layer0_outputs(698)) or (layer0_outputs(6121));
    layer1_outputs(911) <= layer0_outputs(7153);
    layer1_outputs(912) <= (layer0_outputs(4510)) or (layer0_outputs(4493));
    layer1_outputs(913) <= '0';
    layer1_outputs(914) <= not(layer0_outputs(4296));
    layer1_outputs(915) <= not((layer0_outputs(6482)) or (layer0_outputs(3506)));
    layer1_outputs(916) <= layer0_outputs(7921);
    layer1_outputs(917) <= not(layer0_outputs(2248));
    layer1_outputs(918) <= layer0_outputs(7409);
    layer1_outputs(919) <= not(layer0_outputs(8840));
    layer1_outputs(920) <= not((layer0_outputs(3514)) and (layer0_outputs(6418)));
    layer1_outputs(921) <= not(layer0_outputs(7050)) or (layer0_outputs(287));
    layer1_outputs(922) <= '1';
    layer1_outputs(923) <= (layer0_outputs(4991)) and (layer0_outputs(2477));
    layer1_outputs(924) <= layer0_outputs(4390);
    layer1_outputs(925) <= not(layer0_outputs(4085));
    layer1_outputs(926) <= '1';
    layer1_outputs(927) <= layer0_outputs(3803);
    layer1_outputs(928) <= layer0_outputs(2279);
    layer1_outputs(929) <= not((layer0_outputs(6391)) and (layer0_outputs(7035)));
    layer1_outputs(930) <= not(layer0_outputs(9420));
    layer1_outputs(931) <= layer0_outputs(5442);
    layer1_outputs(932) <= (layer0_outputs(5479)) and not (layer0_outputs(4438));
    layer1_outputs(933) <= not((layer0_outputs(9575)) and (layer0_outputs(4495)));
    layer1_outputs(934) <= not((layer0_outputs(5507)) or (layer0_outputs(4247)));
    layer1_outputs(935) <= not((layer0_outputs(7494)) or (layer0_outputs(1794)));
    layer1_outputs(936) <= not(layer0_outputs(4811));
    layer1_outputs(937) <= not((layer0_outputs(2458)) or (layer0_outputs(4131)));
    layer1_outputs(938) <= (layer0_outputs(6103)) and not (layer0_outputs(615));
    layer1_outputs(939) <= not((layer0_outputs(1914)) xor (layer0_outputs(7117)));
    layer1_outputs(940) <= not(layer0_outputs(1589));
    layer1_outputs(941) <= layer0_outputs(3393);
    layer1_outputs(942) <= not(layer0_outputs(4770));
    layer1_outputs(943) <= not((layer0_outputs(5263)) xor (layer0_outputs(9287)));
    layer1_outputs(944) <= not(layer0_outputs(5407));
    layer1_outputs(945) <= layer0_outputs(8691);
    layer1_outputs(946) <= (layer0_outputs(4487)) xor (layer0_outputs(10022));
    layer1_outputs(947) <= (layer0_outputs(10135)) xor (layer0_outputs(1816));
    layer1_outputs(948) <= not(layer0_outputs(7477)) or (layer0_outputs(4429));
    layer1_outputs(949) <= layer0_outputs(1905);
    layer1_outputs(950) <= not(layer0_outputs(6563));
    layer1_outputs(951) <= (layer0_outputs(1216)) and not (layer0_outputs(5691));
    layer1_outputs(952) <= not((layer0_outputs(7758)) and (layer0_outputs(2394)));
    layer1_outputs(953) <= (layer0_outputs(9889)) and not (layer0_outputs(9295));
    layer1_outputs(954) <= (layer0_outputs(8683)) xor (layer0_outputs(1974));
    layer1_outputs(955) <= not((layer0_outputs(6338)) and (layer0_outputs(1850)));
    layer1_outputs(956) <= not(layer0_outputs(3586));
    layer1_outputs(957) <= (layer0_outputs(5321)) or (layer0_outputs(67));
    layer1_outputs(958) <= not(layer0_outputs(2135));
    layer1_outputs(959) <= (layer0_outputs(5419)) and not (layer0_outputs(552));
    layer1_outputs(960) <= (layer0_outputs(947)) and not (layer0_outputs(7742));
    layer1_outputs(961) <= (layer0_outputs(7378)) and (layer0_outputs(10136));
    layer1_outputs(962) <= not(layer0_outputs(2158));
    layer1_outputs(963) <= layer0_outputs(4774);
    layer1_outputs(964) <= layer0_outputs(3600);
    layer1_outputs(965) <= layer0_outputs(5650);
    layer1_outputs(966) <= (layer0_outputs(7843)) xor (layer0_outputs(3790));
    layer1_outputs(967) <= (layer0_outputs(4796)) or (layer0_outputs(4508));
    layer1_outputs(968) <= layer0_outputs(9743);
    layer1_outputs(969) <= not(layer0_outputs(3177)) or (layer0_outputs(5455));
    layer1_outputs(970) <= (layer0_outputs(3716)) and not (layer0_outputs(1491));
    layer1_outputs(971) <= (layer0_outputs(5640)) or (layer0_outputs(2517));
    layer1_outputs(972) <= (layer0_outputs(2610)) and (layer0_outputs(5834));
    layer1_outputs(973) <= '1';
    layer1_outputs(974) <= not((layer0_outputs(9206)) xor (layer0_outputs(8672)));
    layer1_outputs(975) <= layer0_outputs(9767);
    layer1_outputs(976) <= layer0_outputs(7475);
    layer1_outputs(977) <= not(layer0_outputs(4201));
    layer1_outputs(978) <= layer0_outputs(4250);
    layer1_outputs(979) <= (layer0_outputs(184)) and (layer0_outputs(6524));
    layer1_outputs(980) <= not(layer0_outputs(2077));
    layer1_outputs(981) <= layer0_outputs(5372);
    layer1_outputs(982) <= not(layer0_outputs(6522));
    layer1_outputs(983) <= not(layer0_outputs(7998));
    layer1_outputs(984) <= layer0_outputs(9654);
    layer1_outputs(985) <= layer0_outputs(7303);
    layer1_outputs(986) <= not((layer0_outputs(8790)) xor (layer0_outputs(6974)));
    layer1_outputs(987) <= not((layer0_outputs(6923)) and (layer0_outputs(6308)));
    layer1_outputs(988) <= not((layer0_outputs(9015)) and (layer0_outputs(2252)));
    layer1_outputs(989) <= not(layer0_outputs(6004)) or (layer0_outputs(3351));
    layer1_outputs(990) <= layer0_outputs(5578);
    layer1_outputs(991) <= not(layer0_outputs(5352)) or (layer0_outputs(6454));
    layer1_outputs(992) <= layer0_outputs(1507);
    layer1_outputs(993) <= (layer0_outputs(1117)) or (layer0_outputs(7272));
    layer1_outputs(994) <= (layer0_outputs(1464)) and not (layer0_outputs(9189));
    layer1_outputs(995) <= (layer0_outputs(3045)) xor (layer0_outputs(3262));
    layer1_outputs(996) <= (layer0_outputs(1817)) and not (layer0_outputs(915));
    layer1_outputs(997) <= not((layer0_outputs(6068)) and (layer0_outputs(7162)));
    layer1_outputs(998) <= not(layer0_outputs(6840)) or (layer0_outputs(2423));
    layer1_outputs(999) <= (layer0_outputs(6005)) and not (layer0_outputs(3990));
    layer1_outputs(1000) <= not(layer0_outputs(6404));
    layer1_outputs(1001) <= not(layer0_outputs(1853)) or (layer0_outputs(10221));
    layer1_outputs(1002) <= (layer0_outputs(4875)) and not (layer0_outputs(9430));
    layer1_outputs(1003) <= (layer0_outputs(1216)) and not (layer0_outputs(7528));
    layer1_outputs(1004) <= not(layer0_outputs(9612)) or (layer0_outputs(4060));
    layer1_outputs(1005) <= not((layer0_outputs(2274)) or (layer0_outputs(3195)));
    layer1_outputs(1006) <= (layer0_outputs(4436)) and not (layer0_outputs(4087));
    layer1_outputs(1007) <= layer0_outputs(4962);
    layer1_outputs(1008) <= (layer0_outputs(5872)) and not (layer0_outputs(1819));
    layer1_outputs(1009) <= not((layer0_outputs(9620)) and (layer0_outputs(8805)));
    layer1_outputs(1010) <= '1';
    layer1_outputs(1011) <= not(layer0_outputs(3491));
    layer1_outputs(1012) <= not(layer0_outputs(8477)) or (layer0_outputs(8162));
    layer1_outputs(1013) <= (layer0_outputs(2352)) and not (layer0_outputs(978));
    layer1_outputs(1014) <= not(layer0_outputs(4729)) or (layer0_outputs(9912));
    layer1_outputs(1015) <= not(layer0_outputs(7903));
    layer1_outputs(1016) <= not(layer0_outputs(9414));
    layer1_outputs(1017) <= (layer0_outputs(6474)) and (layer0_outputs(4499));
    layer1_outputs(1018) <= not(layer0_outputs(5474));
    layer1_outputs(1019) <= not(layer0_outputs(10172));
    layer1_outputs(1020) <= not(layer0_outputs(10077));
    layer1_outputs(1021) <= (layer0_outputs(6289)) xor (layer0_outputs(9285));
    layer1_outputs(1022) <= not(layer0_outputs(9131));
    layer1_outputs(1023) <= (layer0_outputs(613)) and not (layer0_outputs(3025));
    layer1_outputs(1024) <= not((layer0_outputs(8811)) or (layer0_outputs(1039)));
    layer1_outputs(1025) <= (layer0_outputs(8277)) or (layer0_outputs(1457));
    layer1_outputs(1026) <= not((layer0_outputs(5182)) xor (layer0_outputs(7114)));
    layer1_outputs(1027) <= not(layer0_outputs(3726));
    layer1_outputs(1028) <= '0';
    layer1_outputs(1029) <= (layer0_outputs(5245)) and not (layer0_outputs(1296));
    layer1_outputs(1030) <= not(layer0_outputs(135)) or (layer0_outputs(1192));
    layer1_outputs(1031) <= not((layer0_outputs(4859)) xor (layer0_outputs(8444)));
    layer1_outputs(1032) <= layer0_outputs(7679);
    layer1_outputs(1033) <= not(layer0_outputs(8618)) or (layer0_outputs(8769));
    layer1_outputs(1034) <= not(layer0_outputs(2233)) or (layer0_outputs(7600));
    layer1_outputs(1035) <= (layer0_outputs(2984)) xor (layer0_outputs(4658));
    layer1_outputs(1036) <= (layer0_outputs(5973)) or (layer0_outputs(5858));
    layer1_outputs(1037) <= (layer0_outputs(8462)) and not (layer0_outputs(9510));
    layer1_outputs(1038) <= not(layer0_outputs(4863)) or (layer0_outputs(9863));
    layer1_outputs(1039) <= (layer0_outputs(9234)) and not (layer0_outputs(7022));
    layer1_outputs(1040) <= (layer0_outputs(4946)) xor (layer0_outputs(9365));
    layer1_outputs(1041) <= not((layer0_outputs(5770)) and (layer0_outputs(8514)));
    layer1_outputs(1042) <= (layer0_outputs(4820)) or (layer0_outputs(7350));
    layer1_outputs(1043) <= '0';
    layer1_outputs(1044) <= not(layer0_outputs(3910));
    layer1_outputs(1045) <= (layer0_outputs(6805)) or (layer0_outputs(3676));
    layer1_outputs(1046) <= not(layer0_outputs(10005));
    layer1_outputs(1047) <= (layer0_outputs(9142)) and (layer0_outputs(4681));
    layer1_outputs(1048) <= not(layer0_outputs(1638));
    layer1_outputs(1049) <= layer0_outputs(9356);
    layer1_outputs(1050) <= not((layer0_outputs(5105)) xor (layer0_outputs(1809)));
    layer1_outputs(1051) <= layer0_outputs(8947);
    layer1_outputs(1052) <= not(layer0_outputs(9336));
    layer1_outputs(1053) <= layer0_outputs(3614);
    layer1_outputs(1054) <= not((layer0_outputs(4825)) xor (layer0_outputs(7667)));
    layer1_outputs(1055) <= layer0_outputs(8438);
    layer1_outputs(1056) <= '1';
    layer1_outputs(1057) <= (layer0_outputs(1313)) and not (layer0_outputs(5288));
    layer1_outputs(1058) <= not(layer0_outputs(6039));
    layer1_outputs(1059) <= not(layer0_outputs(6413)) or (layer0_outputs(9139));
    layer1_outputs(1060) <= not(layer0_outputs(7601));
    layer1_outputs(1061) <= (layer0_outputs(6760)) and (layer0_outputs(6789));
    layer1_outputs(1062) <= (layer0_outputs(2786)) or (layer0_outputs(3732));
    layer1_outputs(1063) <= (layer0_outputs(2869)) and not (layer0_outputs(2310));
    layer1_outputs(1064) <= (layer0_outputs(1849)) and not (layer0_outputs(2482));
    layer1_outputs(1065) <= not((layer0_outputs(7576)) and (layer0_outputs(1321)));
    layer1_outputs(1066) <= layer0_outputs(910);
    layer1_outputs(1067) <= not(layer0_outputs(715)) or (layer0_outputs(2493));
    layer1_outputs(1068) <= layer0_outputs(6698);
    layer1_outputs(1069) <= not(layer0_outputs(8766));
    layer1_outputs(1070) <= layer0_outputs(6937);
    layer1_outputs(1071) <= not(layer0_outputs(396));
    layer1_outputs(1072) <= layer0_outputs(2909);
    layer1_outputs(1073) <= (layer0_outputs(1213)) and (layer0_outputs(7098));
    layer1_outputs(1074) <= (layer0_outputs(494)) or (layer0_outputs(3652));
    layer1_outputs(1075) <= not((layer0_outputs(2602)) or (layer0_outputs(8959)));
    layer1_outputs(1076) <= not(layer0_outputs(712)) or (layer0_outputs(1468));
    layer1_outputs(1077) <= not((layer0_outputs(1552)) or (layer0_outputs(8267)));
    layer1_outputs(1078) <= not((layer0_outputs(5374)) xor (layer0_outputs(5031)));
    layer1_outputs(1079) <= layer0_outputs(9325);
    layer1_outputs(1080) <= not(layer0_outputs(4269));
    layer1_outputs(1081) <= layer0_outputs(6411);
    layer1_outputs(1082) <= not(layer0_outputs(6926));
    layer1_outputs(1083) <= '1';
    layer1_outputs(1084) <= not(layer0_outputs(5897));
    layer1_outputs(1085) <= layer0_outputs(10074);
    layer1_outputs(1086) <= not(layer0_outputs(1991));
    layer1_outputs(1087) <= not(layer0_outputs(10163));
    layer1_outputs(1088) <= (layer0_outputs(1110)) or (layer0_outputs(9163));
    layer1_outputs(1089) <= (layer0_outputs(8626)) xor (layer0_outputs(8547));
    layer1_outputs(1090) <= (layer0_outputs(7039)) and not (layer0_outputs(3547));
    layer1_outputs(1091) <= not(layer0_outputs(9291));
    layer1_outputs(1092) <= (layer0_outputs(3926)) and not (layer0_outputs(1768));
    layer1_outputs(1093) <= not((layer0_outputs(7644)) xor (layer0_outputs(5669)));
    layer1_outputs(1094) <= layer0_outputs(4469);
    layer1_outputs(1095) <= not(layer0_outputs(85));
    layer1_outputs(1096) <= not(layer0_outputs(6980));
    layer1_outputs(1097) <= not((layer0_outputs(7280)) or (layer0_outputs(302)));
    layer1_outputs(1098) <= not((layer0_outputs(9262)) or (layer0_outputs(9009)));
    layer1_outputs(1099) <= '1';
    layer1_outputs(1100) <= not((layer0_outputs(4777)) xor (layer0_outputs(9263)));
    layer1_outputs(1101) <= layer0_outputs(4937);
    layer1_outputs(1102) <= not((layer0_outputs(7072)) xor (layer0_outputs(4559)));
    layer1_outputs(1103) <= layer0_outputs(6333);
    layer1_outputs(1104) <= not(layer0_outputs(7640));
    layer1_outputs(1105) <= not(layer0_outputs(8260));
    layer1_outputs(1106) <= layer0_outputs(5537);
    layer1_outputs(1107) <= (layer0_outputs(2384)) and not (layer0_outputs(873));
    layer1_outputs(1108) <= layer0_outputs(3111);
    layer1_outputs(1109) <= layer0_outputs(9594);
    layer1_outputs(1110) <= layer0_outputs(7393);
    layer1_outputs(1111) <= (layer0_outputs(9781)) and not (layer0_outputs(8391));
    layer1_outputs(1112) <= layer0_outputs(8532);
    layer1_outputs(1113) <= not((layer0_outputs(4690)) xor (layer0_outputs(8609)));
    layer1_outputs(1114) <= '1';
    layer1_outputs(1115) <= not((layer0_outputs(6089)) and (layer0_outputs(9919)));
    layer1_outputs(1116) <= not(layer0_outputs(7173)) or (layer0_outputs(5617));
    layer1_outputs(1117) <= not(layer0_outputs(8598));
    layer1_outputs(1118) <= not(layer0_outputs(9574)) or (layer0_outputs(9179));
    layer1_outputs(1119) <= layer0_outputs(4259);
    layer1_outputs(1120) <= '1';
    layer1_outputs(1121) <= (layer0_outputs(771)) and (layer0_outputs(638));
    layer1_outputs(1122) <= (layer0_outputs(6106)) xor (layer0_outputs(5692));
    layer1_outputs(1123) <= (layer0_outputs(1472)) or (layer0_outputs(1339));
    layer1_outputs(1124) <= not((layer0_outputs(9909)) or (layer0_outputs(9792)));
    layer1_outputs(1125) <= not(layer0_outputs(8855)) or (layer0_outputs(8892));
    layer1_outputs(1126) <= not(layer0_outputs(8631));
    layer1_outputs(1127) <= (layer0_outputs(2490)) xor (layer0_outputs(1754));
    layer1_outputs(1128) <= layer0_outputs(8463);
    layer1_outputs(1129) <= layer0_outputs(2453);
    layer1_outputs(1130) <= layer0_outputs(1152);
    layer1_outputs(1131) <= not(layer0_outputs(2511)) or (layer0_outputs(8543));
    layer1_outputs(1132) <= layer0_outputs(7613);
    layer1_outputs(1133) <= (layer0_outputs(3782)) and not (layer0_outputs(2449));
    layer1_outputs(1134) <= layer0_outputs(8217);
    layer1_outputs(1135) <= layer0_outputs(772);
    layer1_outputs(1136) <= not((layer0_outputs(7571)) xor (layer0_outputs(5127)));
    layer1_outputs(1137) <= not(layer0_outputs(9305));
    layer1_outputs(1138) <= layer0_outputs(4599);
    layer1_outputs(1139) <= not(layer0_outputs(2265));
    layer1_outputs(1140) <= not(layer0_outputs(2580)) or (layer0_outputs(9719));
    layer1_outputs(1141) <= (layer0_outputs(2812)) and (layer0_outputs(6438));
    layer1_outputs(1142) <= not(layer0_outputs(8099)) or (layer0_outputs(4699));
    layer1_outputs(1143) <= '1';
    layer1_outputs(1144) <= not(layer0_outputs(8898));
    layer1_outputs(1145) <= not(layer0_outputs(9351));
    layer1_outputs(1146) <= not(layer0_outputs(7273)) or (layer0_outputs(2631));
    layer1_outputs(1147) <= not((layer0_outputs(4050)) or (layer0_outputs(7931)));
    layer1_outputs(1148) <= not((layer0_outputs(6716)) and (layer0_outputs(794)));
    layer1_outputs(1149) <= (layer0_outputs(5271)) and (layer0_outputs(7357));
    layer1_outputs(1150) <= layer0_outputs(8586);
    layer1_outputs(1151) <= (layer0_outputs(9875)) and not (layer0_outputs(1252));
    layer1_outputs(1152) <= not(layer0_outputs(3500)) or (layer0_outputs(8849));
    layer1_outputs(1153) <= not((layer0_outputs(2521)) xor (layer0_outputs(9184)));
    layer1_outputs(1154) <= not(layer0_outputs(8802));
    layer1_outputs(1155) <= (layer0_outputs(6117)) and not (layer0_outputs(9999));
    layer1_outputs(1156) <= layer0_outputs(7157);
    layer1_outputs(1157) <= (layer0_outputs(8901)) and not (layer0_outputs(7099));
    layer1_outputs(1158) <= (layer0_outputs(3544)) and (layer0_outputs(1356));
    layer1_outputs(1159) <= (layer0_outputs(7829)) and not (layer0_outputs(10030));
    layer1_outputs(1160) <= (layer0_outputs(695)) xor (layer0_outputs(7010));
    layer1_outputs(1161) <= layer0_outputs(1087);
    layer1_outputs(1162) <= layer0_outputs(4904);
    layer1_outputs(1163) <= layer0_outputs(9221);
    layer1_outputs(1164) <= (layer0_outputs(435)) or (layer0_outputs(3561));
    layer1_outputs(1165) <= layer0_outputs(3018);
    layer1_outputs(1166) <= not((layer0_outputs(881)) and (layer0_outputs(231)));
    layer1_outputs(1167) <= not((layer0_outputs(457)) and (layer0_outputs(3922)));
    layer1_outputs(1168) <= (layer0_outputs(2956)) and not (layer0_outputs(1088));
    layer1_outputs(1169) <= not((layer0_outputs(10080)) and (layer0_outputs(5899)));
    layer1_outputs(1170) <= '1';
    layer1_outputs(1171) <= not((layer0_outputs(9549)) or (layer0_outputs(9654)));
    layer1_outputs(1172) <= not(layer0_outputs(6776)) or (layer0_outputs(5207));
    layer1_outputs(1173) <= not(layer0_outputs(7571));
    layer1_outputs(1174) <= not(layer0_outputs(2532)) or (layer0_outputs(5141));
    layer1_outputs(1175) <= not(layer0_outputs(5325));
    layer1_outputs(1176) <= not((layer0_outputs(7824)) xor (layer0_outputs(7275)));
    layer1_outputs(1177) <= (layer0_outputs(2512)) and not (layer0_outputs(2888));
    layer1_outputs(1178) <= not((layer0_outputs(4239)) or (layer0_outputs(6729)));
    layer1_outputs(1179) <= not(layer0_outputs(2576)) or (layer0_outputs(8622));
    layer1_outputs(1180) <= (layer0_outputs(3949)) or (layer0_outputs(7567));
    layer1_outputs(1181) <= layer0_outputs(9316);
    layer1_outputs(1182) <= layer0_outputs(4497);
    layer1_outputs(1183) <= (layer0_outputs(9521)) and not (layer0_outputs(9133));
    layer1_outputs(1184) <= not(layer0_outputs(2069)) or (layer0_outputs(6639));
    layer1_outputs(1185) <= (layer0_outputs(7956)) or (layer0_outputs(3728));
    layer1_outputs(1186) <= (layer0_outputs(5104)) and not (layer0_outputs(4777));
    layer1_outputs(1187) <= (layer0_outputs(672)) xor (layer0_outputs(4498));
    layer1_outputs(1188) <= (layer0_outputs(6733)) and not (layer0_outputs(9497));
    layer1_outputs(1189) <= not((layer0_outputs(4261)) and (layer0_outputs(5896)));
    layer1_outputs(1190) <= layer0_outputs(824);
    layer1_outputs(1191) <= not(layer0_outputs(5150)) or (layer0_outputs(9088));
    layer1_outputs(1192) <= layer0_outputs(2891);
    layer1_outputs(1193) <= (layer0_outputs(1842)) and (layer0_outputs(4763));
    layer1_outputs(1194) <= not((layer0_outputs(4522)) or (layer0_outputs(4960)));
    layer1_outputs(1195) <= not(layer0_outputs(9576));
    layer1_outputs(1196) <= layer0_outputs(1263);
    layer1_outputs(1197) <= not((layer0_outputs(6955)) or (layer0_outputs(872)));
    layer1_outputs(1198) <= (layer0_outputs(7165)) and not (layer0_outputs(10233));
    layer1_outputs(1199) <= not(layer0_outputs(9388)) or (layer0_outputs(9257));
    layer1_outputs(1200) <= (layer0_outputs(5713)) xor (layer0_outputs(7827));
    layer1_outputs(1201) <= not(layer0_outputs(8865));
    layer1_outputs(1202) <= not(layer0_outputs(7266));
    layer1_outputs(1203) <= (layer0_outputs(3614)) and not (layer0_outputs(5907));
    layer1_outputs(1204) <= not(layer0_outputs(4649)) or (layer0_outputs(8635));
    layer1_outputs(1205) <= (layer0_outputs(7791)) and (layer0_outputs(3819));
    layer1_outputs(1206) <= not((layer0_outputs(3620)) or (layer0_outputs(9714)));
    layer1_outputs(1207) <= not(layer0_outputs(8611));
    layer1_outputs(1208) <= not((layer0_outputs(2295)) xor (layer0_outputs(4673)));
    layer1_outputs(1209) <= layer0_outputs(6196);
    layer1_outputs(1210) <= not((layer0_outputs(268)) or (layer0_outputs(6052)));
    layer1_outputs(1211) <= not((layer0_outputs(8065)) and (layer0_outputs(7798)));
    layer1_outputs(1212) <= (layer0_outputs(6499)) and not (layer0_outputs(10012));
    layer1_outputs(1213) <= not(layer0_outputs(5952)) or (layer0_outputs(7896));
    layer1_outputs(1214) <= not((layer0_outputs(2093)) and (layer0_outputs(39)));
    layer1_outputs(1215) <= layer0_outputs(2352);
    layer1_outputs(1216) <= layer0_outputs(5795);
    layer1_outputs(1217) <= layer0_outputs(8650);
    layer1_outputs(1218) <= (layer0_outputs(122)) or (layer0_outputs(7423));
    layer1_outputs(1219) <= layer0_outputs(8095);
    layer1_outputs(1220) <= not(layer0_outputs(2732)) or (layer0_outputs(4647));
    layer1_outputs(1221) <= layer0_outputs(4333);
    layer1_outputs(1222) <= (layer0_outputs(2398)) and (layer0_outputs(8059));
    layer1_outputs(1223) <= (layer0_outputs(4145)) xor (layer0_outputs(818));
    layer1_outputs(1224) <= not(layer0_outputs(4182));
    layer1_outputs(1225) <= (layer0_outputs(2378)) and not (layer0_outputs(8882));
    layer1_outputs(1226) <= not(layer0_outputs(7184));
    layer1_outputs(1227) <= (layer0_outputs(4418)) and (layer0_outputs(5398));
    layer1_outputs(1228) <= not(layer0_outputs(2829)) or (layer0_outputs(146));
    layer1_outputs(1229) <= not(layer0_outputs(9530));
    layer1_outputs(1230) <= not((layer0_outputs(609)) or (layer0_outputs(3971)));
    layer1_outputs(1231) <= not(layer0_outputs(9118));
    layer1_outputs(1232) <= layer0_outputs(3665);
    layer1_outputs(1233) <= layer0_outputs(175);
    layer1_outputs(1234) <= (layer0_outputs(501)) xor (layer0_outputs(9590));
    layer1_outputs(1235) <= (layer0_outputs(6558)) and not (layer0_outputs(8237));
    layer1_outputs(1236) <= (layer0_outputs(1915)) xor (layer0_outputs(2244));
    layer1_outputs(1237) <= not(layer0_outputs(3498)) or (layer0_outputs(1421));
    layer1_outputs(1238) <= not((layer0_outputs(5822)) xor (layer0_outputs(8701)));
    layer1_outputs(1239) <= (layer0_outputs(9738)) xor (layer0_outputs(9141));
    layer1_outputs(1240) <= (layer0_outputs(9531)) and not (layer0_outputs(2997));
    layer1_outputs(1241) <= layer0_outputs(7878);
    layer1_outputs(1242) <= (layer0_outputs(3733)) or (layer0_outputs(1437));
    layer1_outputs(1243) <= not((layer0_outputs(401)) or (layer0_outputs(923)));
    layer1_outputs(1244) <= not((layer0_outputs(9504)) and (layer0_outputs(704)));
    layer1_outputs(1245) <= '0';
    layer1_outputs(1246) <= '1';
    layer1_outputs(1247) <= layer0_outputs(6225);
    layer1_outputs(1248) <= layer0_outputs(4622);
    layer1_outputs(1249) <= layer0_outputs(8310);
    layer1_outputs(1250) <= layer0_outputs(3454);
    layer1_outputs(1251) <= (layer0_outputs(4402)) and not (layer0_outputs(766));
    layer1_outputs(1252) <= not((layer0_outputs(6247)) and (layer0_outputs(4439)));
    layer1_outputs(1253) <= not(layer0_outputs(2315));
    layer1_outputs(1254) <= layer0_outputs(866);
    layer1_outputs(1255) <= (layer0_outputs(4664)) and not (layer0_outputs(20));
    layer1_outputs(1256) <= not(layer0_outputs(3530));
    layer1_outputs(1257) <= layer0_outputs(3023);
    layer1_outputs(1258) <= not(layer0_outputs(10054)) or (layer0_outputs(6622));
    layer1_outputs(1259) <= layer0_outputs(7836);
    layer1_outputs(1260) <= (layer0_outputs(9710)) or (layer0_outputs(5289));
    layer1_outputs(1261) <= (layer0_outputs(8243)) or (layer0_outputs(6789));
    layer1_outputs(1262) <= (layer0_outputs(6387)) and (layer0_outputs(5873));
    layer1_outputs(1263) <= not(layer0_outputs(32));
    layer1_outputs(1264) <= (layer0_outputs(4289)) xor (layer0_outputs(8054));
    layer1_outputs(1265) <= (layer0_outputs(2393)) and not (layer0_outputs(971));
    layer1_outputs(1266) <= layer0_outputs(8183);
    layer1_outputs(1267) <= not(layer0_outputs(6647));
    layer1_outputs(1268) <= not((layer0_outputs(4793)) or (layer0_outputs(4069)));
    layer1_outputs(1269) <= layer0_outputs(7629);
    layer1_outputs(1270) <= not(layer0_outputs(3702)) or (layer0_outputs(2763));
    layer1_outputs(1271) <= layer0_outputs(5576);
    layer1_outputs(1272) <= not((layer0_outputs(9035)) and (layer0_outputs(3069)));
    layer1_outputs(1273) <= layer0_outputs(4731);
    layer1_outputs(1274) <= not(layer0_outputs(8734)) or (layer0_outputs(9051));
    layer1_outputs(1275) <= not(layer0_outputs(5367)) or (layer0_outputs(977));
    layer1_outputs(1276) <= (layer0_outputs(3528)) and not (layer0_outputs(2522));
    layer1_outputs(1277) <= not(layer0_outputs(9679));
    layer1_outputs(1278) <= not((layer0_outputs(3753)) or (layer0_outputs(748)));
    layer1_outputs(1279) <= (layer0_outputs(1661)) xor (layer0_outputs(2776));
    layer1_outputs(1280) <= (layer0_outputs(9381)) or (layer0_outputs(3363));
    layer1_outputs(1281) <= not(layer0_outputs(5124));
    layer1_outputs(1282) <= '0';
    layer1_outputs(1283) <= not(layer0_outputs(7435));
    layer1_outputs(1284) <= not(layer0_outputs(4286)) or (layer0_outputs(8455));
    layer1_outputs(1285) <= (layer0_outputs(7370)) and not (layer0_outputs(7894));
    layer1_outputs(1286) <= not(layer0_outputs(7892)) or (layer0_outputs(5565));
    layer1_outputs(1287) <= layer0_outputs(5071);
    layer1_outputs(1288) <= not(layer0_outputs(9399)) or (layer0_outputs(586));
    layer1_outputs(1289) <= (layer0_outputs(4498)) or (layer0_outputs(3577));
    layer1_outputs(1290) <= layer0_outputs(8212);
    layer1_outputs(1291) <= (layer0_outputs(9453)) and not (layer0_outputs(3751));
    layer1_outputs(1292) <= not((layer0_outputs(3511)) or (layer0_outputs(8992)));
    layer1_outputs(1293) <= layer0_outputs(9254);
    layer1_outputs(1294) <= (layer0_outputs(5318)) and (layer0_outputs(3263));
    layer1_outputs(1295) <= not(layer0_outputs(5799));
    layer1_outputs(1296) <= (layer0_outputs(8808)) and not (layer0_outputs(2517));
    layer1_outputs(1297) <= (layer0_outputs(2707)) and not (layer0_outputs(6480));
    layer1_outputs(1298) <= (layer0_outputs(5155)) or (layer0_outputs(10219));
    layer1_outputs(1299) <= (layer0_outputs(3151)) or (layer0_outputs(4153));
    layer1_outputs(1300) <= not(layer0_outputs(2484));
    layer1_outputs(1301) <= not(layer0_outputs(1918)) or (layer0_outputs(9304));
    layer1_outputs(1302) <= (layer0_outputs(4319)) and not (layer0_outputs(4808));
    layer1_outputs(1303) <= not(layer0_outputs(4387));
    layer1_outputs(1304) <= layer0_outputs(2503);
    layer1_outputs(1305) <= (layer0_outputs(4480)) or (layer0_outputs(6753));
    layer1_outputs(1306) <= layer0_outputs(7865);
    layer1_outputs(1307) <= (layer0_outputs(6552)) and (layer0_outputs(4826));
    layer1_outputs(1308) <= not((layer0_outputs(9114)) or (layer0_outputs(4689)));
    layer1_outputs(1309) <= not(layer0_outputs(9547)) or (layer0_outputs(709));
    layer1_outputs(1310) <= (layer0_outputs(5852)) and not (layer0_outputs(7148));
    layer1_outputs(1311) <= not(layer0_outputs(3690));
    layer1_outputs(1312) <= (layer0_outputs(5151)) and not (layer0_outputs(4602));
    layer1_outputs(1313) <= layer0_outputs(7916);
    layer1_outputs(1314) <= (layer0_outputs(2620)) and not (layer0_outputs(7699));
    layer1_outputs(1315) <= layer0_outputs(3325);
    layer1_outputs(1316) <= not((layer0_outputs(8905)) and (layer0_outputs(6191)));
    layer1_outputs(1317) <= (layer0_outputs(7219)) and not (layer0_outputs(7648));
    layer1_outputs(1318) <= layer0_outputs(299);
    layer1_outputs(1319) <= (layer0_outputs(2281)) and not (layer0_outputs(4359));
    layer1_outputs(1320) <= '0';
    layer1_outputs(1321) <= layer0_outputs(5059);
    layer1_outputs(1322) <= layer0_outputs(4445);
    layer1_outputs(1323) <= not(layer0_outputs(7081));
    layer1_outputs(1324) <= not(layer0_outputs(1675));
    layer1_outputs(1325) <= not(layer0_outputs(5485));
    layer1_outputs(1326) <= not((layer0_outputs(923)) and (layer0_outputs(8533)));
    layer1_outputs(1327) <= (layer0_outputs(9721)) and not (layer0_outputs(1600));
    layer1_outputs(1328) <= (layer0_outputs(698)) xor (layer0_outputs(2945));
    layer1_outputs(1329) <= layer0_outputs(4838);
    layer1_outputs(1330) <= not((layer0_outputs(9695)) or (layer0_outputs(7158)));
    layer1_outputs(1331) <= not((layer0_outputs(9917)) and (layer0_outputs(6009)));
    layer1_outputs(1332) <= layer0_outputs(2039);
    layer1_outputs(1333) <= (layer0_outputs(4931)) or (layer0_outputs(1722));
    layer1_outputs(1334) <= (layer0_outputs(5536)) and not (layer0_outputs(4096));
    layer1_outputs(1335) <= not(layer0_outputs(2881));
    layer1_outputs(1336) <= (layer0_outputs(5240)) or (layer0_outputs(8449));
    layer1_outputs(1337) <= (layer0_outputs(5189)) and (layer0_outputs(8972));
    layer1_outputs(1338) <= not((layer0_outputs(7902)) or (layer0_outputs(2465)));
    layer1_outputs(1339) <= layer0_outputs(6646);
    layer1_outputs(1340) <= (layer0_outputs(3518)) and not (layer0_outputs(7317));
    layer1_outputs(1341) <= not((layer0_outputs(2424)) or (layer0_outputs(5745)));
    layer1_outputs(1342) <= (layer0_outputs(1831)) and not (layer0_outputs(4562));
    layer1_outputs(1343) <= layer0_outputs(6793);
    layer1_outputs(1344) <= not((layer0_outputs(1241)) xor (layer0_outputs(2254)));
    layer1_outputs(1345) <= (layer0_outputs(3301)) and not (layer0_outputs(4329));
    layer1_outputs(1346) <= layer0_outputs(2964);
    layer1_outputs(1347) <= not((layer0_outputs(8023)) or (layer0_outputs(3353)));
    layer1_outputs(1348) <= layer0_outputs(7834);
    layer1_outputs(1349) <= not(layer0_outputs(6675)) or (layer0_outputs(8840));
    layer1_outputs(1350) <= not(layer0_outputs(5793)) or (layer0_outputs(2538));
    layer1_outputs(1351) <= not(layer0_outputs(2877)) or (layer0_outputs(7180));
    layer1_outputs(1352) <= layer0_outputs(7566);
    layer1_outputs(1353) <= (layer0_outputs(3974)) and (layer0_outputs(2693));
    layer1_outputs(1354) <= layer0_outputs(5242);
    layer1_outputs(1355) <= layer0_outputs(4064);
    layer1_outputs(1356) <= not(layer0_outputs(7561));
    layer1_outputs(1357) <= (layer0_outputs(2014)) and not (layer0_outputs(453));
    layer1_outputs(1358) <= layer0_outputs(9913);
    layer1_outputs(1359) <= not(layer0_outputs(424)) or (layer0_outputs(3174));
    layer1_outputs(1360) <= not(layer0_outputs(7508)) or (layer0_outputs(8080));
    layer1_outputs(1361) <= layer0_outputs(6772);
    layer1_outputs(1362) <= '0';
    layer1_outputs(1363) <= '0';
    layer1_outputs(1364) <= layer0_outputs(3632);
    layer1_outputs(1365) <= not(layer0_outputs(553)) or (layer0_outputs(3175));
    layer1_outputs(1366) <= not(layer0_outputs(7522)) or (layer0_outputs(7090));
    layer1_outputs(1367) <= not(layer0_outputs(6511)) or (layer0_outputs(3194));
    layer1_outputs(1368) <= layer0_outputs(252);
    layer1_outputs(1369) <= not(layer0_outputs(1953));
    layer1_outputs(1370) <= not(layer0_outputs(2215));
    layer1_outputs(1371) <= not((layer0_outputs(2156)) or (layer0_outputs(8414)));
    layer1_outputs(1372) <= not((layer0_outputs(1063)) or (layer0_outputs(9163)));
    layer1_outputs(1373) <= '1';
    layer1_outputs(1374) <= layer0_outputs(10145);
    layer1_outputs(1375) <= layer0_outputs(8111);
    layer1_outputs(1376) <= '0';
    layer1_outputs(1377) <= not((layer0_outputs(3923)) xor (layer0_outputs(4873)));
    layer1_outputs(1378) <= (layer0_outputs(3464)) or (layer0_outputs(8549));
    layer1_outputs(1379) <= not(layer0_outputs(7044)) or (layer0_outputs(10232));
    layer1_outputs(1380) <= (layer0_outputs(7085)) and not (layer0_outputs(5016));
    layer1_outputs(1381) <= (layer0_outputs(66)) and not (layer0_outputs(464));
    layer1_outputs(1382) <= not(layer0_outputs(267));
    layer1_outputs(1383) <= layer0_outputs(3960);
    layer1_outputs(1384) <= not((layer0_outputs(2330)) xor (layer0_outputs(4900)));
    layer1_outputs(1385) <= not(layer0_outputs(569)) or (layer0_outputs(452));
    layer1_outputs(1386) <= not(layer0_outputs(7513)) or (layer0_outputs(5197));
    layer1_outputs(1387) <= layer0_outputs(9177);
    layer1_outputs(1388) <= (layer0_outputs(685)) and not (layer0_outputs(250));
    layer1_outputs(1389) <= (layer0_outputs(6351)) and not (layer0_outputs(6883));
    layer1_outputs(1390) <= not((layer0_outputs(6453)) or (layer0_outputs(5821)));
    layer1_outputs(1391) <= not(layer0_outputs(6973));
    layer1_outputs(1392) <= not(layer0_outputs(5364));
    layer1_outputs(1393) <= not((layer0_outputs(2260)) or (layer0_outputs(7723)));
    layer1_outputs(1394) <= (layer0_outputs(7321)) or (layer0_outputs(6608));
    layer1_outputs(1395) <= not(layer0_outputs(10099));
    layer1_outputs(1396) <= not(layer0_outputs(341)) or (layer0_outputs(5059));
    layer1_outputs(1397) <= not(layer0_outputs(4799)) or (layer0_outputs(3048));
    layer1_outputs(1398) <= '0';
    layer1_outputs(1399) <= (layer0_outputs(9036)) and not (layer0_outputs(8599));
    layer1_outputs(1400) <= (layer0_outputs(4119)) xor (layer0_outputs(7321));
    layer1_outputs(1401) <= not((layer0_outputs(4901)) xor (layer0_outputs(6286)));
    layer1_outputs(1402) <= layer0_outputs(8085);
    layer1_outputs(1403) <= not((layer0_outputs(2725)) xor (layer0_outputs(10235)));
    layer1_outputs(1404) <= not((layer0_outputs(1812)) or (layer0_outputs(4741)));
    layer1_outputs(1405) <= (layer0_outputs(8761)) and not (layer0_outputs(6995));
    layer1_outputs(1406) <= layer0_outputs(8231);
    layer1_outputs(1407) <= not((layer0_outputs(5530)) xor (layer0_outputs(8316)));
    layer1_outputs(1408) <= layer0_outputs(1656);
    layer1_outputs(1409) <= layer0_outputs(4188);
    layer1_outputs(1410) <= not(layer0_outputs(4607)) or (layer0_outputs(576));
    layer1_outputs(1411) <= not(layer0_outputs(6812));
    layer1_outputs(1412) <= not((layer0_outputs(4629)) xor (layer0_outputs(9741)));
    layer1_outputs(1413) <= not(layer0_outputs(2116));
    layer1_outputs(1414) <= not(layer0_outputs(4812));
    layer1_outputs(1415) <= not(layer0_outputs(4377));
    layer1_outputs(1416) <= (layer0_outputs(6649)) and not (layer0_outputs(7964));
    layer1_outputs(1417) <= (layer0_outputs(5515)) xor (layer0_outputs(4855));
    layer1_outputs(1418) <= not(layer0_outputs(2328));
    layer1_outputs(1419) <= not((layer0_outputs(1891)) and (layer0_outputs(1648)));
    layer1_outputs(1420) <= not((layer0_outputs(8450)) or (layer0_outputs(2160)));
    layer1_outputs(1421) <= not(layer0_outputs(8042));
    layer1_outputs(1422) <= not(layer0_outputs(9815));
    layer1_outputs(1423) <= layer0_outputs(5849);
    layer1_outputs(1424) <= not(layer0_outputs(8213)) or (layer0_outputs(6625));
    layer1_outputs(1425) <= '1';
    layer1_outputs(1426) <= (layer0_outputs(3854)) or (layer0_outputs(2063));
    layer1_outputs(1427) <= (layer0_outputs(8541)) or (layer0_outputs(2526));
    layer1_outputs(1428) <= not(layer0_outputs(6986)) or (layer0_outputs(1649));
    layer1_outputs(1429) <= layer0_outputs(8493);
    layer1_outputs(1430) <= '1';
    layer1_outputs(1431) <= '0';
    layer1_outputs(1432) <= not(layer0_outputs(6313)) or (layer0_outputs(6710));
    layer1_outputs(1433) <= not((layer0_outputs(9344)) xor (layer0_outputs(1903)));
    layer1_outputs(1434) <= not((layer0_outputs(6303)) xor (layer0_outputs(9941)));
    layer1_outputs(1435) <= (layer0_outputs(9899)) and not (layer0_outputs(248));
    layer1_outputs(1436) <= not((layer0_outputs(1858)) xor (layer0_outputs(29)));
    layer1_outputs(1437) <= '0';
    layer1_outputs(1438) <= not(layer0_outputs(4202)) or (layer0_outputs(87));
    layer1_outputs(1439) <= not(layer0_outputs(1569)) or (layer0_outputs(8793));
    layer1_outputs(1440) <= not((layer0_outputs(5033)) or (layer0_outputs(613)));
    layer1_outputs(1441) <= layer0_outputs(580);
    layer1_outputs(1442) <= not((layer0_outputs(2917)) and (layer0_outputs(10079)));
    layer1_outputs(1443) <= not((layer0_outputs(6111)) and (layer0_outputs(6711)));
    layer1_outputs(1444) <= (layer0_outputs(501)) or (layer0_outputs(381));
    layer1_outputs(1445) <= not((layer0_outputs(5350)) or (layer0_outputs(5329)));
    layer1_outputs(1446) <= not(layer0_outputs(3616)) or (layer0_outputs(4506));
    layer1_outputs(1447) <= (layer0_outputs(5234)) and not (layer0_outputs(7138));
    layer1_outputs(1448) <= (layer0_outputs(1310)) and not (layer0_outputs(1911));
    layer1_outputs(1449) <= not(layer0_outputs(1147));
    layer1_outputs(1450) <= layer0_outputs(4042);
    layer1_outputs(1451) <= not((layer0_outputs(5874)) and (layer0_outputs(2060)));
    layer1_outputs(1452) <= layer0_outputs(7299);
    layer1_outputs(1453) <= (layer0_outputs(1207)) or (layer0_outputs(7291));
    layer1_outputs(1454) <= not(layer0_outputs(8659));
    layer1_outputs(1455) <= not((layer0_outputs(2356)) xor (layer0_outputs(8377)));
    layer1_outputs(1456) <= not(layer0_outputs(5208));
    layer1_outputs(1457) <= layer0_outputs(288);
    layer1_outputs(1458) <= layer0_outputs(7018);
    layer1_outputs(1459) <= (layer0_outputs(2322)) and (layer0_outputs(8126));
    layer1_outputs(1460) <= layer0_outputs(1437);
    layer1_outputs(1461) <= (layer0_outputs(2679)) xor (layer0_outputs(2249));
    layer1_outputs(1462) <= (layer0_outputs(178)) and not (layer0_outputs(7001));
    layer1_outputs(1463) <= layer0_outputs(372);
    layer1_outputs(1464) <= not((layer0_outputs(6403)) or (layer0_outputs(7921)));
    layer1_outputs(1465) <= (layer0_outputs(2526)) and not (layer0_outputs(4082));
    layer1_outputs(1466) <= layer0_outputs(8251);
    layer1_outputs(1467) <= not(layer0_outputs(9300));
    layer1_outputs(1468) <= not(layer0_outputs(6748)) or (layer0_outputs(4100));
    layer1_outputs(1469) <= not((layer0_outputs(7397)) xor (layer0_outputs(5975)));
    layer1_outputs(1470) <= not(layer0_outputs(8864)) or (layer0_outputs(412));
    layer1_outputs(1471) <= layer0_outputs(8736);
    layer1_outputs(1472) <= not((layer0_outputs(4633)) and (layer0_outputs(1574)));
    layer1_outputs(1473) <= not(layer0_outputs(404)) or (layer0_outputs(7163));
    layer1_outputs(1474) <= (layer0_outputs(9201)) or (layer0_outputs(3616));
    layer1_outputs(1475) <= (layer0_outputs(9167)) and (layer0_outputs(7278));
    layer1_outputs(1476) <= (layer0_outputs(5614)) and not (layer0_outputs(5399));
    layer1_outputs(1477) <= layer0_outputs(4637);
    layer1_outputs(1478) <= layer0_outputs(4726);
    layer1_outputs(1479) <= (layer0_outputs(6267)) and not (layer0_outputs(1593));
    layer1_outputs(1480) <= (layer0_outputs(9617)) and not (layer0_outputs(98));
    layer1_outputs(1481) <= not(layer0_outputs(4779));
    layer1_outputs(1482) <= (layer0_outputs(2860)) and not (layer0_outputs(3373));
    layer1_outputs(1483) <= (layer0_outputs(1824)) or (layer0_outputs(8554));
    layer1_outputs(1484) <= not(layer0_outputs(10016));
    layer1_outputs(1485) <= (layer0_outputs(9078)) and (layer0_outputs(6710));
    layer1_outputs(1486) <= (layer0_outputs(9495)) or (layer0_outputs(1499));
    layer1_outputs(1487) <= (layer0_outputs(701)) or (layer0_outputs(8797));
    layer1_outputs(1488) <= not(layer0_outputs(5951));
    layer1_outputs(1489) <= not((layer0_outputs(9565)) and (layer0_outputs(2073)));
    layer1_outputs(1490) <= (layer0_outputs(8813)) and not (layer0_outputs(9383));
    layer1_outputs(1491) <= (layer0_outputs(1325)) or (layer0_outputs(9764));
    layer1_outputs(1492) <= (layer0_outputs(7413)) xor (layer0_outputs(9088));
    layer1_outputs(1493) <= layer0_outputs(2337);
    layer1_outputs(1494) <= not(layer0_outputs(3022));
    layer1_outputs(1495) <= not(layer0_outputs(9259));
    layer1_outputs(1496) <= not(layer0_outputs(1460));
    layer1_outputs(1497) <= (layer0_outputs(8868)) and not (layer0_outputs(1651));
    layer1_outputs(1498) <= '1';
    layer1_outputs(1499) <= not(layer0_outputs(9280)) or (layer0_outputs(9497));
    layer1_outputs(1500) <= not((layer0_outputs(5310)) or (layer0_outputs(8549)));
    layer1_outputs(1501) <= not((layer0_outputs(6021)) xor (layer0_outputs(3701)));
    layer1_outputs(1502) <= layer0_outputs(7276);
    layer1_outputs(1503) <= not(layer0_outputs(9210));
    layer1_outputs(1504) <= layer0_outputs(6413);
    layer1_outputs(1505) <= (layer0_outputs(7088)) and not (layer0_outputs(6075));
    layer1_outputs(1506) <= not(layer0_outputs(8027));
    layer1_outputs(1507) <= not(layer0_outputs(4205)) or (layer0_outputs(3561));
    layer1_outputs(1508) <= not((layer0_outputs(9104)) or (layer0_outputs(4273)));
    layer1_outputs(1509) <= (layer0_outputs(941)) and not (layer0_outputs(5323));
    layer1_outputs(1510) <= (layer0_outputs(1932)) and (layer0_outputs(1578));
    layer1_outputs(1511) <= (layer0_outputs(8425)) and not (layer0_outputs(2191));
    layer1_outputs(1512) <= not(layer0_outputs(7213)) or (layer0_outputs(8521));
    layer1_outputs(1513) <= (layer0_outputs(2305)) and not (layer0_outputs(4120));
    layer1_outputs(1514) <= layer0_outputs(9854);
    layer1_outputs(1515) <= (layer0_outputs(2093)) and (layer0_outputs(1792));
    layer1_outputs(1516) <= not((layer0_outputs(4910)) xor (layer0_outputs(3285)));
    layer1_outputs(1517) <= not(layer0_outputs(9147));
    layer1_outputs(1518) <= (layer0_outputs(4883)) or (layer0_outputs(2456));
    layer1_outputs(1519) <= not(layer0_outputs(10036));
    layer1_outputs(1520) <= not((layer0_outputs(2341)) or (layer0_outputs(7652)));
    layer1_outputs(1521) <= not((layer0_outputs(6587)) and (layer0_outputs(1310)));
    layer1_outputs(1522) <= not(layer0_outputs(8980));
    layer1_outputs(1523) <= not(layer0_outputs(7575));
    layer1_outputs(1524) <= not(layer0_outputs(3715)) or (layer0_outputs(2316));
    layer1_outputs(1525) <= (layer0_outputs(632)) and not (layer0_outputs(7287));
    layer1_outputs(1526) <= not((layer0_outputs(8583)) xor (layer0_outputs(6963)));
    layer1_outputs(1527) <= not(layer0_outputs(2081));
    layer1_outputs(1528) <= (layer0_outputs(9328)) or (layer0_outputs(390));
    layer1_outputs(1529) <= not(layer0_outputs(3298)) or (layer0_outputs(6326));
    layer1_outputs(1530) <= not(layer0_outputs(5663));
    layer1_outputs(1531) <= layer0_outputs(10027);
    layer1_outputs(1532) <= layer0_outputs(1005);
    layer1_outputs(1533) <= not(layer0_outputs(1480));
    layer1_outputs(1534) <= not((layer0_outputs(1161)) and (layer0_outputs(5107)));
    layer1_outputs(1535) <= (layer0_outputs(5804)) or (layer0_outputs(3847));
    layer1_outputs(1536) <= not(layer0_outputs(8553));
    layer1_outputs(1537) <= (layer0_outputs(1484)) and (layer0_outputs(6578));
    layer1_outputs(1538) <= not(layer0_outputs(8319));
    layer1_outputs(1539) <= not((layer0_outputs(1768)) or (layer0_outputs(8902)));
    layer1_outputs(1540) <= not(layer0_outputs(1254));
    layer1_outputs(1541) <= not(layer0_outputs(4099));
    layer1_outputs(1542) <= not((layer0_outputs(6982)) xor (layer0_outputs(4326)));
    layer1_outputs(1543) <= (layer0_outputs(8437)) or (layer0_outputs(5025));
    layer1_outputs(1544) <= not(layer0_outputs(218)) or (layer0_outputs(8527));
    layer1_outputs(1545) <= not(layer0_outputs(2400)) or (layer0_outputs(7146));
    layer1_outputs(1546) <= '0';
    layer1_outputs(1547) <= layer0_outputs(3304);
    layer1_outputs(1548) <= (layer0_outputs(1287)) and (layer0_outputs(10147));
    layer1_outputs(1549) <= not(layer0_outputs(5160));
    layer1_outputs(1550) <= not(layer0_outputs(1367));
    layer1_outputs(1551) <= (layer0_outputs(3379)) and not (layer0_outputs(5295));
    layer1_outputs(1552) <= not(layer0_outputs(10237));
    layer1_outputs(1553) <= not(layer0_outputs(8392));
    layer1_outputs(1554) <= (layer0_outputs(3305)) xor (layer0_outputs(3981));
    layer1_outputs(1555) <= (layer0_outputs(6543)) or (layer0_outputs(1110));
    layer1_outputs(1556) <= (layer0_outputs(8386)) and not (layer0_outputs(9577));
    layer1_outputs(1557) <= not(layer0_outputs(6212));
    layer1_outputs(1558) <= not((layer0_outputs(5941)) and (layer0_outputs(5369)));
    layer1_outputs(1559) <= not(layer0_outputs(2585)) or (layer0_outputs(1297));
    layer1_outputs(1560) <= not(layer0_outputs(9319));
    layer1_outputs(1561) <= not(layer0_outputs(9217));
    layer1_outputs(1562) <= layer0_outputs(4598);
    layer1_outputs(1563) <= not((layer0_outputs(6499)) xor (layer0_outputs(7426)));
    layer1_outputs(1564) <= not(layer0_outputs(1640));
    layer1_outputs(1565) <= layer0_outputs(9537);
    layer1_outputs(1566) <= not(layer0_outputs(8494));
    layer1_outputs(1567) <= not(layer0_outputs(6578));
    layer1_outputs(1568) <= '0';
    layer1_outputs(1569) <= not((layer0_outputs(5888)) and (layer0_outputs(873)));
    layer1_outputs(1570) <= not(layer0_outputs(8922));
    layer1_outputs(1571) <= not(layer0_outputs(10003));
    layer1_outputs(1572) <= (layer0_outputs(5689)) xor (layer0_outputs(808));
    layer1_outputs(1573) <= layer0_outputs(9573);
    layer1_outputs(1574) <= not(layer0_outputs(1556)) or (layer0_outputs(3295));
    layer1_outputs(1575) <= not(layer0_outputs(5166)) or (layer0_outputs(1394));
    layer1_outputs(1576) <= not(layer0_outputs(3276));
    layer1_outputs(1577) <= not((layer0_outputs(2486)) or (layer0_outputs(463)));
    layer1_outputs(1578) <= (layer0_outputs(1541)) xor (layer0_outputs(895));
    layer1_outputs(1579) <= (layer0_outputs(3128)) and not (layer0_outputs(7048));
    layer1_outputs(1580) <= '0';
    layer1_outputs(1581) <= '1';
    layer1_outputs(1582) <= not(layer0_outputs(4939));
    layer1_outputs(1583) <= not((layer0_outputs(659)) and (layer0_outputs(7922)));
    layer1_outputs(1584) <= layer0_outputs(4286);
    layer1_outputs(1585) <= '0';
    layer1_outputs(1586) <= not(layer0_outputs(3940));
    layer1_outputs(1587) <= not((layer0_outputs(458)) xor (layer0_outputs(8441)));
    layer1_outputs(1588) <= layer0_outputs(3899);
    layer1_outputs(1589) <= layer0_outputs(3036);
    layer1_outputs(1590) <= (layer0_outputs(4386)) or (layer0_outputs(1323));
    layer1_outputs(1591) <= not((layer0_outputs(4189)) or (layer0_outputs(2626)));
    layer1_outputs(1592) <= not(layer0_outputs(147));
    layer1_outputs(1593) <= layer0_outputs(834);
    layer1_outputs(1594) <= (layer0_outputs(7871)) or (layer0_outputs(7237));
    layer1_outputs(1595) <= not(layer0_outputs(4539));
    layer1_outputs(1596) <= not(layer0_outputs(7346));
    layer1_outputs(1597) <= (layer0_outputs(5083)) and not (layer0_outputs(1993));
    layer1_outputs(1598) <= not(layer0_outputs(1667));
    layer1_outputs(1599) <= not(layer0_outputs(2414)) or (layer0_outputs(8050));
    layer1_outputs(1600) <= (layer0_outputs(9219)) and (layer0_outputs(1111));
    layer1_outputs(1601) <= (layer0_outputs(6215)) and (layer0_outputs(8452));
    layer1_outputs(1602) <= not((layer0_outputs(4348)) or (layer0_outputs(6894)));
    layer1_outputs(1603) <= (layer0_outputs(3399)) and not (layer0_outputs(3743));
    layer1_outputs(1604) <= not(layer0_outputs(5630));
    layer1_outputs(1605) <= not((layer0_outputs(4376)) or (layer0_outputs(4336)));
    layer1_outputs(1606) <= not(layer0_outputs(1467)) or (layer0_outputs(807));
    layer1_outputs(1607) <= not((layer0_outputs(2260)) and (layer0_outputs(2960)));
    layer1_outputs(1608) <= not(layer0_outputs(6152));
    layer1_outputs(1609) <= not(layer0_outputs(2231));
    layer1_outputs(1610) <= not(layer0_outputs(3403));
    layer1_outputs(1611) <= layer0_outputs(6372);
    layer1_outputs(1612) <= not(layer0_outputs(5743));
    layer1_outputs(1613) <= not(layer0_outputs(5378));
    layer1_outputs(1614) <= '0';
    layer1_outputs(1615) <= '0';
    layer1_outputs(1616) <= (layer0_outputs(7383)) and (layer0_outputs(8546));
    layer1_outputs(1617) <= (layer0_outputs(5034)) and not (layer0_outputs(5670));
    layer1_outputs(1618) <= (layer0_outputs(415)) xor (layer0_outputs(9609));
    layer1_outputs(1619) <= (layer0_outputs(3278)) or (layer0_outputs(6666));
    layer1_outputs(1620) <= not(layer0_outputs(3450));
    layer1_outputs(1621) <= not((layer0_outputs(2381)) xor (layer0_outputs(6447)));
    layer1_outputs(1622) <= (layer0_outputs(5728)) and not (layer0_outputs(3772));
    layer1_outputs(1623) <= layer0_outputs(8231);
    layer1_outputs(1624) <= not((layer0_outputs(1031)) or (layer0_outputs(2785)));
    layer1_outputs(1625) <= layer0_outputs(1183);
    layer1_outputs(1626) <= not(layer0_outputs(4526));
    layer1_outputs(1627) <= not((layer0_outputs(4896)) and (layer0_outputs(6265)));
    layer1_outputs(1628) <= (layer0_outputs(1460)) and (layer0_outputs(1314));
    layer1_outputs(1629) <= not((layer0_outputs(4021)) or (layer0_outputs(8054)));
    layer1_outputs(1630) <= (layer0_outputs(2198)) or (layer0_outputs(2070));
    layer1_outputs(1631) <= not(layer0_outputs(8604)) or (layer0_outputs(5506));
    layer1_outputs(1632) <= not(layer0_outputs(8694));
    layer1_outputs(1633) <= not((layer0_outputs(1282)) or (layer0_outputs(7923)));
    layer1_outputs(1634) <= '0';
    layer1_outputs(1635) <= (layer0_outputs(819)) and (layer0_outputs(101));
    layer1_outputs(1636) <= not(layer0_outputs(8182));
    layer1_outputs(1637) <= not((layer0_outputs(7243)) xor (layer0_outputs(199)));
    layer1_outputs(1638) <= (layer0_outputs(8408)) and not (layer0_outputs(2571));
    layer1_outputs(1639) <= not(layer0_outputs(3163));
    layer1_outputs(1640) <= (layer0_outputs(5779)) and (layer0_outputs(9447));
    layer1_outputs(1641) <= not(layer0_outputs(7601));
    layer1_outputs(1642) <= (layer0_outputs(950)) and not (layer0_outputs(5676));
    layer1_outputs(1643) <= (layer0_outputs(243)) and not (layer0_outputs(3045));
    layer1_outputs(1644) <= (layer0_outputs(8296)) and not (layer0_outputs(1760));
    layer1_outputs(1645) <= not(layer0_outputs(567));
    layer1_outputs(1646) <= layer0_outputs(1039);
    layer1_outputs(1647) <= (layer0_outputs(7968)) and not (layer0_outputs(1416));
    layer1_outputs(1648) <= layer0_outputs(8867);
    layer1_outputs(1649) <= layer0_outputs(2853);
    layer1_outputs(1650) <= (layer0_outputs(9242)) and not (layer0_outputs(3411));
    layer1_outputs(1651) <= (layer0_outputs(8176)) and (layer0_outputs(9775));
    layer1_outputs(1652) <= (layer0_outputs(7803)) and not (layer0_outputs(6659));
    layer1_outputs(1653) <= not((layer0_outputs(7599)) and (layer0_outputs(10067)));
    layer1_outputs(1654) <= not(layer0_outputs(589));
    layer1_outputs(1655) <= not((layer0_outputs(7581)) xor (layer0_outputs(2892)));
    layer1_outputs(1656) <= layer0_outputs(1619);
    layer1_outputs(1657) <= not(layer0_outputs(6137));
    layer1_outputs(1658) <= (layer0_outputs(4895)) xor (layer0_outputs(8582));
    layer1_outputs(1659) <= not(layer0_outputs(6082));
    layer1_outputs(1660) <= (layer0_outputs(8711)) and not (layer0_outputs(8876));
    layer1_outputs(1661) <= (layer0_outputs(581)) and not (layer0_outputs(392));
    layer1_outputs(1662) <= not((layer0_outputs(1134)) and (layer0_outputs(1194)));
    layer1_outputs(1663) <= layer0_outputs(9290);
    layer1_outputs(1664) <= '1';
    layer1_outputs(1665) <= layer0_outputs(5655);
    layer1_outputs(1666) <= layer0_outputs(2719);
    layer1_outputs(1667) <= not(layer0_outputs(4483)) or (layer0_outputs(1230));
    layer1_outputs(1668) <= layer0_outputs(4970);
    layer1_outputs(1669) <= (layer0_outputs(6656)) and not (layer0_outputs(4226));
    layer1_outputs(1670) <= (layer0_outputs(3484)) xor (layer0_outputs(2342));
    layer1_outputs(1671) <= layer0_outputs(4735);
    layer1_outputs(1672) <= not((layer0_outputs(4530)) or (layer0_outputs(7623)));
    layer1_outputs(1673) <= (layer0_outputs(515)) xor (layer0_outputs(10014));
    layer1_outputs(1674) <= not((layer0_outputs(1975)) xor (layer0_outputs(814)));
    layer1_outputs(1675) <= (layer0_outputs(8851)) and (layer0_outputs(7522));
    layer1_outputs(1676) <= not((layer0_outputs(4213)) xor (layer0_outputs(4076)));
    layer1_outputs(1677) <= layer0_outputs(4596);
    layer1_outputs(1678) <= not(layer0_outputs(4646));
    layer1_outputs(1679) <= '1';
    layer1_outputs(1680) <= (layer0_outputs(9774)) and not (layer0_outputs(646));
    layer1_outputs(1681) <= layer0_outputs(710);
    layer1_outputs(1682) <= not(layer0_outputs(528));
    layer1_outputs(1683) <= not(layer0_outputs(6209)) or (layer0_outputs(8358));
    layer1_outputs(1684) <= not(layer0_outputs(8669)) or (layer0_outputs(9819));
    layer1_outputs(1685) <= layer0_outputs(5725);
    layer1_outputs(1686) <= layer0_outputs(9108);
    layer1_outputs(1687) <= layer0_outputs(2494);
    layer1_outputs(1688) <= not(layer0_outputs(1912)) or (layer0_outputs(2801));
    layer1_outputs(1689) <= layer0_outputs(5094);
    layer1_outputs(1690) <= layer0_outputs(1720);
    layer1_outputs(1691) <= not((layer0_outputs(4625)) and (layer0_outputs(8103)));
    layer1_outputs(1692) <= not(layer0_outputs(4418));
    layer1_outputs(1693) <= not(layer0_outputs(1833));
    layer1_outputs(1694) <= not((layer0_outputs(8817)) xor (layer0_outputs(9600)));
    layer1_outputs(1695) <= not(layer0_outputs(2085));
    layer1_outputs(1696) <= not(layer0_outputs(5712));
    layer1_outputs(1697) <= not(layer0_outputs(3089)) or (layer0_outputs(1916));
    layer1_outputs(1698) <= not(layer0_outputs(8582));
    layer1_outputs(1699) <= (layer0_outputs(8062)) and not (layer0_outputs(9587));
    layer1_outputs(1700) <= not(layer0_outputs(1027));
    layer1_outputs(1701) <= (layer0_outputs(1900)) and not (layer0_outputs(6023));
    layer1_outputs(1702) <= (layer0_outputs(6324)) and not (layer0_outputs(5005));
    layer1_outputs(1703) <= not(layer0_outputs(2210)) or (layer0_outputs(1345));
    layer1_outputs(1704) <= (layer0_outputs(9627)) or (layer0_outputs(2761));
    layer1_outputs(1705) <= not((layer0_outputs(2199)) xor (layer0_outputs(9842)));
    layer1_outputs(1706) <= layer0_outputs(2968);
    layer1_outputs(1707) <= (layer0_outputs(6267)) and not (layer0_outputs(4050));
    layer1_outputs(1708) <= (layer0_outputs(2638)) or (layer0_outputs(2404));
    layer1_outputs(1709) <= not((layer0_outputs(4375)) and (layer0_outputs(8259)));
    layer1_outputs(1710) <= not((layer0_outputs(1247)) xor (layer0_outputs(1452)));
    layer1_outputs(1711) <= not(layer0_outputs(6076));
    layer1_outputs(1712) <= not(layer0_outputs(7979));
    layer1_outputs(1713) <= layer0_outputs(5880);
    layer1_outputs(1714) <= (layer0_outputs(1031)) or (layer0_outputs(7455));
    layer1_outputs(1715) <= '0';
    layer1_outputs(1716) <= not(layer0_outputs(7196));
    layer1_outputs(1717) <= layer0_outputs(10210);
    layer1_outputs(1718) <= not(layer0_outputs(5355));
    layer1_outputs(1719) <= (layer0_outputs(6813)) xor (layer0_outputs(9300));
    layer1_outputs(1720) <= not(layer0_outputs(9525));
    layer1_outputs(1721) <= not(layer0_outputs(5810));
    layer1_outputs(1722) <= not(layer0_outputs(784));
    layer1_outputs(1723) <= layer0_outputs(7778);
    layer1_outputs(1724) <= not(layer0_outputs(320));
    layer1_outputs(1725) <= (layer0_outputs(3073)) and not (layer0_outputs(706));
    layer1_outputs(1726) <= not(layer0_outputs(36)) or (layer0_outputs(9859));
    layer1_outputs(1727) <= not(layer0_outputs(7335)) or (layer0_outputs(3799));
    layer1_outputs(1728) <= (layer0_outputs(1690)) and (layer0_outputs(4950));
    layer1_outputs(1729) <= not((layer0_outputs(3570)) or (layer0_outputs(6834)));
    layer1_outputs(1730) <= not(layer0_outputs(6365));
    layer1_outputs(1731) <= not(layer0_outputs(1225));
    layer1_outputs(1732) <= (layer0_outputs(7189)) or (layer0_outputs(3099));
    layer1_outputs(1733) <= layer0_outputs(7789);
    layer1_outputs(1734) <= not(layer0_outputs(1244));
    layer1_outputs(1735) <= not(layer0_outputs(5014));
    layer1_outputs(1736) <= (layer0_outputs(2803)) and not (layer0_outputs(4954));
    layer1_outputs(1737) <= layer0_outputs(8015);
    layer1_outputs(1738) <= layer0_outputs(7773);
    layer1_outputs(1739) <= (layer0_outputs(942)) xor (layer0_outputs(5531));
    layer1_outputs(1740) <= (layer0_outputs(2870)) and not (layer0_outputs(2119));
    layer1_outputs(1741) <= not(layer0_outputs(908));
    layer1_outputs(1742) <= not(layer0_outputs(7241));
    layer1_outputs(1743) <= not(layer0_outputs(9424)) or (layer0_outputs(9396));
    layer1_outputs(1744) <= (layer0_outputs(5520)) and not (layer0_outputs(5069));
    layer1_outputs(1745) <= (layer0_outputs(10041)) and (layer0_outputs(7453));
    layer1_outputs(1746) <= not(layer0_outputs(9203)) or (layer0_outputs(2009));
    layer1_outputs(1747) <= not(layer0_outputs(7352));
    layer1_outputs(1748) <= (layer0_outputs(8029)) and (layer0_outputs(2099));
    layer1_outputs(1749) <= (layer0_outputs(6679)) or (layer0_outputs(7779));
    layer1_outputs(1750) <= layer0_outputs(6525);
    layer1_outputs(1751) <= not(layer0_outputs(2755));
    layer1_outputs(1752) <= (layer0_outputs(2701)) and not (layer0_outputs(8774));
    layer1_outputs(1753) <= (layer0_outputs(1617)) and not (layer0_outputs(892));
    layer1_outputs(1754) <= (layer0_outputs(7067)) and not (layer0_outputs(3956));
    layer1_outputs(1755) <= not(layer0_outputs(7)) or (layer0_outputs(1339));
    layer1_outputs(1756) <= (layer0_outputs(2955)) or (layer0_outputs(4934));
    layer1_outputs(1757) <= layer0_outputs(8487);
    layer1_outputs(1758) <= layer0_outputs(9578);
    layer1_outputs(1759) <= layer0_outputs(6407);
    layer1_outputs(1760) <= layer0_outputs(7514);
    layer1_outputs(1761) <= not(layer0_outputs(9888));
    layer1_outputs(1762) <= (layer0_outputs(2553)) and (layer0_outputs(3366));
    layer1_outputs(1763) <= layer0_outputs(6744);
    layer1_outputs(1764) <= not(layer0_outputs(6550)) or (layer0_outputs(3043));
    layer1_outputs(1765) <= (layer0_outputs(4947)) or (layer0_outputs(1084));
    layer1_outputs(1766) <= (layer0_outputs(9281)) and not (layer0_outputs(6797));
    layer1_outputs(1767) <= not((layer0_outputs(7169)) or (layer0_outputs(257)));
    layer1_outputs(1768) <= not(layer0_outputs(9197)) or (layer0_outputs(8916));
    layer1_outputs(1769) <= not(layer0_outputs(10200));
    layer1_outputs(1770) <= layer0_outputs(8145);
    layer1_outputs(1771) <= (layer0_outputs(8434)) or (layer0_outputs(3715));
    layer1_outputs(1772) <= (layer0_outputs(541)) xor (layer0_outputs(8371));
    layer1_outputs(1773) <= (layer0_outputs(4854)) xor (layer0_outputs(6410));
    layer1_outputs(1774) <= '1';
    layer1_outputs(1775) <= not((layer0_outputs(3335)) and (layer0_outputs(393)));
    layer1_outputs(1776) <= not(layer0_outputs(9176)) or (layer0_outputs(4210));
    layer1_outputs(1777) <= '0';
    layer1_outputs(1778) <= not(layer0_outputs(804));
    layer1_outputs(1779) <= not(layer0_outputs(1923));
    layer1_outputs(1780) <= not((layer0_outputs(1563)) and (layer0_outputs(2401)));
    layer1_outputs(1781) <= not(layer0_outputs(6637));
    layer1_outputs(1782) <= (layer0_outputs(6490)) and not (layer0_outputs(348));
    layer1_outputs(1783) <= (layer0_outputs(1653)) and (layer0_outputs(9677));
    layer1_outputs(1784) <= not(layer0_outputs(2752)) or (layer0_outputs(7621));
    layer1_outputs(1785) <= not((layer0_outputs(6957)) or (layer0_outputs(2614)));
    layer1_outputs(1786) <= not((layer0_outputs(10018)) or (layer0_outputs(1513)));
    layer1_outputs(1787) <= layer0_outputs(4292);
    layer1_outputs(1788) <= (layer0_outputs(5470)) and not (layer0_outputs(1857));
    layer1_outputs(1789) <= not(layer0_outputs(4255));
    layer1_outputs(1790) <= not(layer0_outputs(1530));
    layer1_outputs(1791) <= layer0_outputs(9646);
    layer1_outputs(1792) <= (layer0_outputs(1820)) and not (layer0_outputs(3456));
    layer1_outputs(1793) <= not((layer0_outputs(2445)) and (layer0_outputs(4277)));
    layer1_outputs(1794) <= not(layer0_outputs(612));
    layer1_outputs(1795) <= layer0_outputs(7660);
    layer1_outputs(1796) <= (layer0_outputs(7787)) and not (layer0_outputs(6010));
    layer1_outputs(1797) <= layer0_outputs(4426);
    layer1_outputs(1798) <= not(layer0_outputs(6299));
    layer1_outputs(1799) <= not(layer0_outputs(8435));
    layer1_outputs(1800) <= not(layer0_outputs(4738)) or (layer0_outputs(9650));
    layer1_outputs(1801) <= not(layer0_outputs(8527));
    layer1_outputs(1802) <= not(layer0_outputs(5596));
    layer1_outputs(1803) <= not(layer0_outputs(3434)) or (layer0_outputs(6909));
    layer1_outputs(1804) <= (layer0_outputs(2930)) and not (layer0_outputs(4774));
    layer1_outputs(1805) <= not((layer0_outputs(3965)) and (layer0_outputs(4804)));
    layer1_outputs(1806) <= not((layer0_outputs(10139)) or (layer0_outputs(550)));
    layer1_outputs(1807) <= not(layer0_outputs(8593));
    layer1_outputs(1808) <= not((layer0_outputs(5747)) or (layer0_outputs(946)));
    layer1_outputs(1809) <= (layer0_outputs(6691)) xor (layer0_outputs(37));
    layer1_outputs(1810) <= not(layer0_outputs(1023));
    layer1_outputs(1811) <= (layer0_outputs(5332)) and not (layer0_outputs(1793));
    layer1_outputs(1812) <= not(layer0_outputs(6198));
    layer1_outputs(1813) <= (layer0_outputs(6174)) and not (layer0_outputs(6021));
    layer1_outputs(1814) <= not(layer0_outputs(5198)) or (layer0_outputs(2153));
    layer1_outputs(1815) <= not((layer0_outputs(888)) or (layer0_outputs(4344)));
    layer1_outputs(1816) <= (layer0_outputs(3257)) xor (layer0_outputs(6161));
    layer1_outputs(1817) <= layer0_outputs(6270);
    layer1_outputs(1818) <= (layer0_outputs(3807)) and (layer0_outputs(5829));
    layer1_outputs(1819) <= layer0_outputs(6496);
    layer1_outputs(1820) <= not(layer0_outputs(6247));
    layer1_outputs(1821) <= (layer0_outputs(408)) or (layer0_outputs(6094));
    layer1_outputs(1822) <= layer0_outputs(10211);
    layer1_outputs(1823) <= layer0_outputs(5064);
    layer1_outputs(1824) <= not(layer0_outputs(1485));
    layer1_outputs(1825) <= not((layer0_outputs(8198)) and (layer0_outputs(2002)));
    layer1_outputs(1826) <= not((layer0_outputs(10051)) and (layer0_outputs(9952)));
    layer1_outputs(1827) <= layer0_outputs(5723);
    layer1_outputs(1828) <= not((layer0_outputs(3106)) or (layer0_outputs(8573)));
    layer1_outputs(1829) <= (layer0_outputs(2620)) and (layer0_outputs(7995));
    layer1_outputs(1830) <= layer0_outputs(3977);
    layer1_outputs(1831) <= (layer0_outputs(4379)) and (layer0_outputs(1482));
    layer1_outputs(1832) <= not((layer0_outputs(6647)) xor (layer0_outputs(2756)));
    layer1_outputs(1833) <= not(layer0_outputs(6775));
    layer1_outputs(1834) <= layer0_outputs(4859);
    layer1_outputs(1835) <= not((layer0_outputs(9750)) xor (layer0_outputs(2172)));
    layer1_outputs(1836) <= not(layer0_outputs(4122));
    layer1_outputs(1837) <= (layer0_outputs(4122)) and (layer0_outputs(2280));
    layer1_outputs(1838) <= layer0_outputs(7785);
    layer1_outputs(1839) <= not(layer0_outputs(4395));
    layer1_outputs(1840) <= not((layer0_outputs(42)) and (layer0_outputs(867)));
    layer1_outputs(1841) <= (layer0_outputs(5020)) and not (layer0_outputs(1796));
    layer1_outputs(1842) <= not(layer0_outputs(7432));
    layer1_outputs(1843) <= layer0_outputs(1586);
    layer1_outputs(1844) <= not(layer0_outputs(8185));
    layer1_outputs(1845) <= not((layer0_outputs(9993)) xor (layer0_outputs(6034)));
    layer1_outputs(1846) <= '1';
    layer1_outputs(1847) <= layer0_outputs(7054);
    layer1_outputs(1848) <= not(layer0_outputs(2714));
    layer1_outputs(1849) <= not(layer0_outputs(5960));
    layer1_outputs(1850) <= (layer0_outputs(4604)) or (layer0_outputs(3193));
    layer1_outputs(1851) <= layer0_outputs(6990);
    layer1_outputs(1852) <= (layer0_outputs(5683)) and (layer0_outputs(1970));
    layer1_outputs(1853) <= (layer0_outputs(5203)) xor (layer0_outputs(775));
    layer1_outputs(1854) <= not(layer0_outputs(2100));
    layer1_outputs(1855) <= (layer0_outputs(5986)) and not (layer0_outputs(4174));
    layer1_outputs(1856) <= not((layer0_outputs(6162)) and (layer0_outputs(10113)));
    layer1_outputs(1857) <= not(layer0_outputs(3407));
    layer1_outputs(1858) <= not((layer0_outputs(6492)) xor (layer0_outputs(5174)));
    layer1_outputs(1859) <= not((layer0_outputs(9488)) and (layer0_outputs(4641)));
    layer1_outputs(1860) <= layer0_outputs(5193);
    layer1_outputs(1861) <= '1';
    layer1_outputs(1862) <= not(layer0_outputs(9156));
    layer1_outputs(1863) <= not((layer0_outputs(8319)) or (layer0_outputs(5313)));
    layer1_outputs(1864) <= not(layer0_outputs(10022)) or (layer0_outputs(5990));
    layer1_outputs(1865) <= not((layer0_outputs(5014)) xor (layer0_outputs(9523)));
    layer1_outputs(1866) <= not(layer0_outputs(6562));
    layer1_outputs(1867) <= (layer0_outputs(7368)) and not (layer0_outputs(1009));
    layer1_outputs(1868) <= layer0_outputs(7093);
    layer1_outputs(1869) <= (layer0_outputs(1293)) and not (layer0_outputs(3312));
    layer1_outputs(1870) <= '1';
    layer1_outputs(1871) <= layer0_outputs(811);
    layer1_outputs(1872) <= (layer0_outputs(6099)) or (layer0_outputs(9796));
    layer1_outputs(1873) <= (layer0_outputs(3129)) and not (layer0_outputs(5672));
    layer1_outputs(1874) <= (layer0_outputs(6586)) or (layer0_outputs(7947));
    layer1_outputs(1875) <= layer0_outputs(4070);
    layer1_outputs(1876) <= not((layer0_outputs(9207)) and (layer0_outputs(3367)));
    layer1_outputs(1877) <= layer0_outputs(7125);
    layer1_outputs(1878) <= (layer0_outputs(5437)) or (layer0_outputs(6246));
    layer1_outputs(1879) <= (layer0_outputs(7970)) and not (layer0_outputs(4524));
    layer1_outputs(1880) <= not((layer0_outputs(4327)) or (layer0_outputs(10123)));
    layer1_outputs(1881) <= (layer0_outputs(191)) and not (layer0_outputs(9284));
    layer1_outputs(1882) <= not(layer0_outputs(4888));
    layer1_outputs(1883) <= not((layer0_outputs(6453)) or (layer0_outputs(2736)));
    layer1_outputs(1884) <= (layer0_outputs(4358)) xor (layer0_outputs(9452));
    layer1_outputs(1885) <= not(layer0_outputs(8897)) or (layer0_outputs(5065));
    layer1_outputs(1886) <= (layer0_outputs(502)) and not (layer0_outputs(6660));
    layer1_outputs(1887) <= not((layer0_outputs(5487)) or (layer0_outputs(6412)));
    layer1_outputs(1888) <= not(layer0_outputs(6885));
    layer1_outputs(1889) <= not(layer0_outputs(1649));
    layer1_outputs(1890) <= (layer0_outputs(3245)) and not (layer0_outputs(7683));
    layer1_outputs(1891) <= not((layer0_outputs(8081)) and (layer0_outputs(1388)));
    layer1_outputs(1892) <= (layer0_outputs(2989)) or (layer0_outputs(7));
    layer1_outputs(1893) <= (layer0_outputs(8285)) and (layer0_outputs(8853));
    layer1_outputs(1894) <= not((layer0_outputs(7957)) xor (layer0_outputs(9620)));
    layer1_outputs(1895) <= not(layer0_outputs(8265)) or (layer0_outputs(6202));
    layer1_outputs(1896) <= not(layer0_outputs(6414));
    layer1_outputs(1897) <= not(layer0_outputs(1367));
    layer1_outputs(1898) <= not(layer0_outputs(4207));
    layer1_outputs(1899) <= layer0_outputs(1289);
    layer1_outputs(1900) <= layer0_outputs(858);
    layer1_outputs(1901) <= (layer0_outputs(2715)) or (layer0_outputs(7706));
    layer1_outputs(1902) <= (layer0_outputs(6567)) and not (layer0_outputs(9533));
    layer1_outputs(1903) <= layer0_outputs(4768);
    layer1_outputs(1904) <= layer0_outputs(3727);
    layer1_outputs(1905) <= (layer0_outputs(5085)) or (layer0_outputs(3305));
    layer1_outputs(1906) <= (layer0_outputs(295)) and (layer0_outputs(9466));
    layer1_outputs(1907) <= (layer0_outputs(10209)) and not (layer0_outputs(2985));
    layer1_outputs(1908) <= layer0_outputs(7294);
    layer1_outputs(1909) <= not(layer0_outputs(2469)) or (layer0_outputs(1813));
    layer1_outputs(1910) <= (layer0_outputs(625)) and (layer0_outputs(554));
    layer1_outputs(1911) <= layer0_outputs(4989);
    layer1_outputs(1912) <= not(layer0_outputs(8567)) or (layer0_outputs(1051));
    layer1_outputs(1913) <= not(layer0_outputs(9411));
    layer1_outputs(1914) <= (layer0_outputs(9864)) and (layer0_outputs(6411));
    layer1_outputs(1915) <= layer0_outputs(3294);
    layer1_outputs(1916) <= (layer0_outputs(8538)) and not (layer0_outputs(5830));
    layer1_outputs(1917) <= layer0_outputs(6838);
    layer1_outputs(1918) <= '1';
    layer1_outputs(1919) <= (layer0_outputs(3898)) or (layer0_outputs(4182));
    layer1_outputs(1920) <= not(layer0_outputs(31));
    layer1_outputs(1921) <= not((layer0_outputs(9476)) and (layer0_outputs(5124)));
    layer1_outputs(1922) <= (layer0_outputs(9623)) xor (layer0_outputs(852));
    layer1_outputs(1923) <= not(layer0_outputs(9));
    layer1_outputs(1924) <= not((layer0_outputs(1596)) xor (layer0_outputs(8879)));
    layer1_outputs(1925) <= (layer0_outputs(6443)) and (layer0_outputs(4283));
    layer1_outputs(1926) <= layer0_outputs(9203);
    layer1_outputs(1927) <= not((layer0_outputs(4861)) and (layer0_outputs(5062)));
    layer1_outputs(1928) <= not((layer0_outputs(5)) xor (layer0_outputs(7478)));
    layer1_outputs(1929) <= not((layer0_outputs(453)) and (layer0_outputs(2918)));
    layer1_outputs(1930) <= not(layer0_outputs(2771));
    layer1_outputs(1931) <= layer0_outputs(8405);
    layer1_outputs(1932) <= layer0_outputs(7060);
    layer1_outputs(1933) <= not(layer0_outputs(8937));
    layer1_outputs(1934) <= (layer0_outputs(6941)) and (layer0_outputs(6842));
    layer1_outputs(1935) <= not(layer0_outputs(5467));
    layer1_outputs(1936) <= not(layer0_outputs(4392));
    layer1_outputs(1937) <= (layer0_outputs(7317)) xor (layer0_outputs(8008));
    layer1_outputs(1938) <= not(layer0_outputs(2061)) or (layer0_outputs(8935));
    layer1_outputs(1939) <= layer0_outputs(2340);
    layer1_outputs(1940) <= not((layer0_outputs(4669)) and (layer0_outputs(608)));
    layer1_outputs(1941) <= '1';
    layer1_outputs(1942) <= (layer0_outputs(3024)) and not (layer0_outputs(7173));
    layer1_outputs(1943) <= not(layer0_outputs(7031));
    layer1_outputs(1944) <= layer0_outputs(9639);
    layer1_outputs(1945) <= not((layer0_outputs(1299)) and (layer0_outputs(8498)));
    layer1_outputs(1946) <= not((layer0_outputs(9438)) or (layer0_outputs(5400)));
    layer1_outputs(1947) <= not(layer0_outputs(6336)) or (layer0_outputs(4913));
    layer1_outputs(1948) <= (layer0_outputs(7328)) or (layer0_outputs(5734));
    layer1_outputs(1949) <= not(layer0_outputs(7853)) or (layer0_outputs(5038));
    layer1_outputs(1950) <= not(layer0_outputs(1447));
    layer1_outputs(1951) <= (layer0_outputs(3608)) and not (layer0_outputs(5832));
    layer1_outputs(1952) <= (layer0_outputs(378)) and not (layer0_outputs(3812));
    layer1_outputs(1953) <= (layer0_outputs(622)) and (layer0_outputs(3168));
    layer1_outputs(1954) <= (layer0_outputs(9154)) and (layer0_outputs(7359));
    layer1_outputs(1955) <= (layer0_outputs(7110)) and not (layer0_outputs(2520));
    layer1_outputs(1956) <= not((layer0_outputs(9524)) and (layer0_outputs(160)));
    layer1_outputs(1957) <= (layer0_outputs(1730)) xor (layer0_outputs(2285));
    layer1_outputs(1958) <= (layer0_outputs(9240)) or (layer0_outputs(649));
    layer1_outputs(1959) <= layer0_outputs(1330);
    layer1_outputs(1960) <= '1';
    layer1_outputs(1961) <= not(layer0_outputs(9759)) or (layer0_outputs(6533));
    layer1_outputs(1962) <= layer0_outputs(8771);
    layer1_outputs(1963) <= (layer0_outputs(5607)) and (layer0_outputs(835));
    layer1_outputs(1964) <= (layer0_outputs(7411)) and not (layer0_outputs(1799));
    layer1_outputs(1965) <= not((layer0_outputs(2108)) and (layer0_outputs(5759)));
    layer1_outputs(1966) <= not(layer0_outputs(2941));
    layer1_outputs(1967) <= layer0_outputs(919);
    layer1_outputs(1968) <= layer0_outputs(121);
    layer1_outputs(1969) <= not((layer0_outputs(1563)) or (layer0_outputs(4492)));
    layer1_outputs(1970) <= not(layer0_outputs(4532)) or (layer0_outputs(8966));
    layer1_outputs(1971) <= not((layer0_outputs(1759)) and (layer0_outputs(5514)));
    layer1_outputs(1972) <= layer0_outputs(6381);
    layer1_outputs(1973) <= not(layer0_outputs(3302)) or (layer0_outputs(7911));
    layer1_outputs(1974) <= not(layer0_outputs(1771));
    layer1_outputs(1975) <= layer0_outputs(30);
    layer1_outputs(1976) <= layer0_outputs(266);
    layer1_outputs(1977) <= not((layer0_outputs(7401)) or (layer0_outputs(3406)));
    layer1_outputs(1978) <= not(layer0_outputs(6208)) or (layer0_outputs(9103));
    layer1_outputs(1979) <= not((layer0_outputs(4490)) xor (layer0_outputs(8809)));
    layer1_outputs(1980) <= not((layer0_outputs(148)) or (layer0_outputs(5769)));
    layer1_outputs(1981) <= not(layer0_outputs(7023)) or (layer0_outputs(4458));
    layer1_outputs(1982) <= (layer0_outputs(619)) and not (layer0_outputs(1035));
    layer1_outputs(1983) <= not(layer0_outputs(5652)) or (layer0_outputs(4259));
    layer1_outputs(1984) <= (layer0_outputs(2428)) and not (layer0_outputs(3759));
    layer1_outputs(1985) <= not(layer0_outputs(8766));
    layer1_outputs(1986) <= not(layer0_outputs(6817));
    layer1_outputs(1987) <= not(layer0_outputs(8574));
    layer1_outputs(1988) <= layer0_outputs(1522);
    layer1_outputs(1989) <= not(layer0_outputs(3472)) or (layer0_outputs(7821));
    layer1_outputs(1990) <= (layer0_outputs(8718)) and not (layer0_outputs(8623));
    layer1_outputs(1991) <= (layer0_outputs(8033)) and not (layer0_outputs(832));
    layer1_outputs(1992) <= not(layer0_outputs(6913));
    layer1_outputs(1993) <= layer0_outputs(9271);
    layer1_outputs(1994) <= not((layer0_outputs(6594)) and (layer0_outputs(2456)));
    layer1_outputs(1995) <= not((layer0_outputs(1353)) and (layer0_outputs(8036)));
    layer1_outputs(1996) <= not((layer0_outputs(5987)) xor (layer0_outputs(9132)));
    layer1_outputs(1997) <= (layer0_outputs(9595)) and not (layer0_outputs(1259));
    layer1_outputs(1998) <= not((layer0_outputs(7471)) or (layer0_outputs(9115)));
    layer1_outputs(1999) <= not(layer0_outputs(1958));
    layer1_outputs(2000) <= not((layer0_outputs(850)) and (layer0_outputs(9629)));
    layer1_outputs(2001) <= layer0_outputs(7040);
    layer1_outputs(2002) <= (layer0_outputs(4929)) or (layer0_outputs(4066));
    layer1_outputs(2003) <= (layer0_outputs(5868)) and (layer0_outputs(2298));
    layer1_outputs(2004) <= layer0_outputs(6175);
    layer1_outputs(2005) <= layer0_outputs(5991);
    layer1_outputs(2006) <= not((layer0_outputs(7470)) or (layer0_outputs(1797)));
    layer1_outputs(2007) <= not(layer0_outputs(3128));
    layer1_outputs(2008) <= (layer0_outputs(9932)) xor (layer0_outputs(10146));
    layer1_outputs(2009) <= not(layer0_outputs(8673));
    layer1_outputs(2010) <= not(layer0_outputs(6203));
    layer1_outputs(2011) <= layer0_outputs(3255);
    layer1_outputs(2012) <= not((layer0_outputs(2378)) and (layer0_outputs(3621)));
    layer1_outputs(2013) <= (layer0_outputs(4532)) and not (layer0_outputs(8843));
    layer1_outputs(2014) <= not((layer0_outputs(5081)) xor (layer0_outputs(8164)));
    layer1_outputs(2015) <= (layer0_outputs(5589)) and (layer0_outputs(290));
    layer1_outputs(2016) <= not(layer0_outputs(1055)) or (layer0_outputs(6046));
    layer1_outputs(2017) <= not((layer0_outputs(5604)) and (layer0_outputs(6753)));
    layer1_outputs(2018) <= (layer0_outputs(9270)) xor (layer0_outputs(4645));
    layer1_outputs(2019) <= (layer0_outputs(10162)) or (layer0_outputs(43));
    layer1_outputs(2020) <= (layer0_outputs(9717)) and not (layer0_outputs(8774));
    layer1_outputs(2021) <= '0';
    layer1_outputs(2022) <= '0';
    layer1_outputs(2023) <= not(layer0_outputs(7954)) or (layer0_outputs(9449));
    layer1_outputs(2024) <= '0';
    layer1_outputs(2025) <= layer0_outputs(6152);
    layer1_outputs(2026) <= not(layer0_outputs(3525));
    layer1_outputs(2027) <= not((layer0_outputs(1163)) and (layer0_outputs(7393)));
    layer1_outputs(2028) <= not((layer0_outputs(4534)) and (layer0_outputs(5252)));
    layer1_outputs(2029) <= layer0_outputs(8049);
    layer1_outputs(2030) <= (layer0_outputs(9046)) and not (layer0_outputs(8359));
    layer1_outputs(2031) <= not(layer0_outputs(5010));
    layer1_outputs(2032) <= (layer0_outputs(8744)) and not (layer0_outputs(5259));
    layer1_outputs(2033) <= not(layer0_outputs(2882));
    layer1_outputs(2034) <= not((layer0_outputs(355)) xor (layer0_outputs(1304)));
    layer1_outputs(2035) <= not(layer0_outputs(1711));
    layer1_outputs(2036) <= not((layer0_outputs(1564)) or (layer0_outputs(8064)));
    layer1_outputs(2037) <= layer0_outputs(3012);
    layer1_outputs(2038) <= (layer0_outputs(6872)) and (layer0_outputs(2387));
    layer1_outputs(2039) <= (layer0_outputs(3755)) xor (layer0_outputs(5401));
    layer1_outputs(2040) <= not(layer0_outputs(8215)) or (layer0_outputs(6464));
    layer1_outputs(2041) <= layer0_outputs(2538);
    layer1_outputs(2042) <= layer0_outputs(2603);
    layer1_outputs(2043) <= not(layer0_outputs(10214));
    layer1_outputs(2044) <= (layer0_outputs(7747)) xor (layer0_outputs(9532));
    layer1_outputs(2045) <= layer0_outputs(4505);
    layer1_outputs(2046) <= layer0_outputs(4002);
    layer1_outputs(2047) <= (layer0_outputs(2)) xor (layer0_outputs(2204));
    layer1_outputs(2048) <= (layer0_outputs(1535)) and (layer0_outputs(5999));
    layer1_outputs(2049) <= not((layer0_outputs(10072)) xor (layer0_outputs(3044)));
    layer1_outputs(2050) <= (layer0_outputs(264)) or (layer0_outputs(9863));
    layer1_outputs(2051) <= layer0_outputs(3087);
    layer1_outputs(2052) <= layer0_outputs(2554);
    layer1_outputs(2053) <= not(layer0_outputs(6069));
    layer1_outputs(2054) <= (layer0_outputs(6444)) or (layer0_outputs(519));
    layer1_outputs(2055) <= not(layer0_outputs(2625));
    layer1_outputs(2056) <= not(layer0_outputs(9728)) or (layer0_outputs(6862));
    layer1_outputs(2057) <= not(layer0_outputs(9269));
    layer1_outputs(2058) <= not(layer0_outputs(9288));
    layer1_outputs(2059) <= (layer0_outputs(8011)) xor (layer0_outputs(6687));
    layer1_outputs(2060) <= (layer0_outputs(7885)) and not (layer0_outputs(1832));
    layer1_outputs(2061) <= not((layer0_outputs(480)) xor (layer0_outputs(4872)));
    layer1_outputs(2062) <= not(layer0_outputs(2327));
    layer1_outputs(2063) <= not(layer0_outputs(2486));
    layer1_outputs(2064) <= not(layer0_outputs(4580)) or (layer0_outputs(9970));
    layer1_outputs(2065) <= (layer0_outputs(5417)) xor (layer0_outputs(6263));
    layer1_outputs(2066) <= (layer0_outputs(5883)) and (layer0_outputs(7192));
    layer1_outputs(2067) <= not(layer0_outputs(6737));
    layer1_outputs(2068) <= not(layer0_outputs(7615));
    layer1_outputs(2069) <= layer0_outputs(9374);
    layer1_outputs(2070) <= layer0_outputs(2790);
    layer1_outputs(2071) <= not((layer0_outputs(8884)) xor (layer0_outputs(9229)));
    layer1_outputs(2072) <= (layer0_outputs(10019)) and (layer0_outputs(8967));
    layer1_outputs(2073) <= '0';
    layer1_outputs(2074) <= (layer0_outputs(9049)) and not (layer0_outputs(949));
    layer1_outputs(2075) <= (layer0_outputs(3189)) and not (layer0_outputs(823));
    layer1_outputs(2076) <= not(layer0_outputs(5301)) or (layer0_outputs(5165));
    layer1_outputs(2077) <= not(layer0_outputs(8214));
    layer1_outputs(2078) <= layer0_outputs(9119);
    layer1_outputs(2079) <= layer0_outputs(10165);
    layer1_outputs(2080) <= layer0_outputs(5857);
    layer1_outputs(2081) <= not((layer0_outputs(6508)) and (layer0_outputs(6151)));
    layer1_outputs(2082) <= not((layer0_outputs(3252)) xor (layer0_outputs(1184)));
    layer1_outputs(2083) <= not(layer0_outputs(1846)) or (layer0_outputs(4661));
    layer1_outputs(2084) <= (layer0_outputs(9933)) and (layer0_outputs(9179));
    layer1_outputs(2085) <= not((layer0_outputs(4351)) and (layer0_outputs(4321)));
    layer1_outputs(2086) <= (layer0_outputs(4097)) xor (layer0_outputs(1682));
    layer1_outputs(2087) <= layer0_outputs(8305);
    layer1_outputs(2088) <= layer0_outputs(3773);
    layer1_outputs(2089) <= not((layer0_outputs(3757)) or (layer0_outputs(26)));
    layer1_outputs(2090) <= not(layer0_outputs(9821));
    layer1_outputs(2091) <= not(layer0_outputs(5903));
    layer1_outputs(2092) <= (layer0_outputs(8042)) and not (layer0_outputs(7293));
    layer1_outputs(2093) <= layer0_outputs(326);
    layer1_outputs(2094) <= not((layer0_outputs(7342)) xor (layer0_outputs(1979)));
    layer1_outputs(2095) <= not(layer0_outputs(8909));
    layer1_outputs(2096) <= not((layer0_outputs(5347)) or (layer0_outputs(3028)));
    layer1_outputs(2097) <= not(layer0_outputs(1067)) or (layer0_outputs(6617));
    layer1_outputs(2098) <= (layer0_outputs(9454)) and not (layer0_outputs(9528));
    layer1_outputs(2099) <= not(layer0_outputs(5870));
    layer1_outputs(2100) <= not((layer0_outputs(5317)) xor (layer0_outputs(5706)));
    layer1_outputs(2101) <= layer0_outputs(137);
    layer1_outputs(2102) <= layer0_outputs(1580);
    layer1_outputs(2103) <= (layer0_outputs(2016)) and not (layer0_outputs(6427));
    layer1_outputs(2104) <= (layer0_outputs(9312)) xor (layer0_outputs(5756));
    layer1_outputs(2105) <= not((layer0_outputs(6500)) and (layer0_outputs(9247)));
    layer1_outputs(2106) <= not(layer0_outputs(5807));
    layer1_outputs(2107) <= not(layer0_outputs(6282));
    layer1_outputs(2108) <= (layer0_outputs(8261)) and (layer0_outputs(2346));
    layer1_outputs(2109) <= layer0_outputs(8010);
    layer1_outputs(2110) <= (layer0_outputs(5926)) xor (layer0_outputs(2651));
    layer1_outputs(2111) <= (layer0_outputs(1802)) and (layer0_outputs(8870));
    layer1_outputs(2112) <= not((layer0_outputs(6884)) xor (layer0_outputs(6502)));
    layer1_outputs(2113) <= layer0_outputs(3668);
    layer1_outputs(2114) <= layer0_outputs(7534);
    layer1_outputs(2115) <= not((layer0_outputs(9878)) and (layer0_outputs(2978)));
    layer1_outputs(2116) <= layer0_outputs(3606);
    layer1_outputs(2117) <= (layer0_outputs(662)) xor (layer0_outputs(4961));
    layer1_outputs(2118) <= not((layer0_outputs(141)) or (layer0_outputs(2245)));
    layer1_outputs(2119) <= (layer0_outputs(6293)) xor (layer0_outputs(3659));
    layer1_outputs(2120) <= not((layer0_outputs(8587)) or (layer0_outputs(4204)));
    layer1_outputs(2121) <= not(layer0_outputs(1785));
    layer1_outputs(2122) <= not(layer0_outputs(8758));
    layer1_outputs(2123) <= (layer0_outputs(878)) and (layer0_outputs(9882));
    layer1_outputs(2124) <= not((layer0_outputs(9089)) xor (layer0_outputs(5458)));
    layer1_outputs(2125) <= (layer0_outputs(2588)) and not (layer0_outputs(8297));
    layer1_outputs(2126) <= not((layer0_outputs(4781)) or (layer0_outputs(4807)));
    layer1_outputs(2127) <= (layer0_outputs(5009)) xor (layer0_outputs(37));
    layer1_outputs(2128) <= layer0_outputs(8347);
    layer1_outputs(2129) <= (layer0_outputs(7416)) and (layer0_outputs(620));
    layer1_outputs(2130) <= not(layer0_outputs(1781)) or (layer0_outputs(1869));
    layer1_outputs(2131) <= (layer0_outputs(7546)) or (layer0_outputs(7469));
    layer1_outputs(2132) <= not(layer0_outputs(3332));
    layer1_outputs(2133) <= layer0_outputs(3681);
    layer1_outputs(2134) <= layer0_outputs(7920);
    layer1_outputs(2135) <= not(layer0_outputs(7287));
    layer1_outputs(2136) <= (layer0_outputs(1929)) and not (layer0_outputs(9631));
    layer1_outputs(2137) <= not(layer0_outputs(2654));
    layer1_outputs(2138) <= layer0_outputs(5703);
    layer1_outputs(2139) <= layer0_outputs(9414);
    layer1_outputs(2140) <= (layer0_outputs(7385)) or (layer0_outputs(2555));
    layer1_outputs(2141) <= (layer0_outputs(6148)) xor (layer0_outputs(820));
    layer1_outputs(2142) <= not(layer0_outputs(9804));
    layer1_outputs(2143) <= (layer0_outputs(3369)) and (layer0_outputs(7611));
    layer1_outputs(2144) <= not((layer0_outputs(562)) and (layer0_outputs(9058)));
    layer1_outputs(2145) <= (layer0_outputs(2036)) and (layer0_outputs(7990));
    layer1_outputs(2146) <= layer0_outputs(8895);
    layer1_outputs(2147) <= not((layer0_outputs(7181)) and (layer0_outputs(10087)));
    layer1_outputs(2148) <= not(layer0_outputs(822));
    layer1_outputs(2149) <= not((layer0_outputs(7568)) xor (layer0_outputs(1160)));
    layer1_outputs(2150) <= not((layer0_outputs(4691)) and (layer0_outputs(786)));
    layer1_outputs(2151) <= layer0_outputs(8764);
    layer1_outputs(2152) <= (layer0_outputs(2117)) and not (layer0_outputs(10154));
    layer1_outputs(2153) <= not(layer0_outputs(8994));
    layer1_outputs(2154) <= not(layer0_outputs(3697));
    layer1_outputs(2155) <= not(layer0_outputs(585));
    layer1_outputs(2156) <= (layer0_outputs(9703)) and (layer0_outputs(6461));
    layer1_outputs(2157) <= not(layer0_outputs(4330));
    layer1_outputs(2158) <= not(layer0_outputs(1173));
    layer1_outputs(2159) <= layer0_outputs(4827);
    layer1_outputs(2160) <= (layer0_outputs(7692)) and not (layer0_outputs(5046));
    layer1_outputs(2161) <= (layer0_outputs(3899)) and not (layer0_outputs(6778));
    layer1_outputs(2162) <= not((layer0_outputs(1791)) and (layer0_outputs(59)));
    layer1_outputs(2163) <= (layer0_outputs(4448)) and not (layer0_outputs(3251));
    layer1_outputs(2164) <= not(layer0_outputs(3656)) or (layer0_outputs(3662));
    layer1_outputs(2165) <= not((layer0_outputs(7577)) or (layer0_outputs(5476)));
    layer1_outputs(2166) <= not((layer0_outputs(8508)) and (layer0_outputs(1316)));
    layer1_outputs(2167) <= not(layer0_outputs(6081)) or (layer0_outputs(9960));
    layer1_outputs(2168) <= (layer0_outputs(5412)) or (layer0_outputs(6820));
    layer1_outputs(2169) <= not(layer0_outputs(712));
    layer1_outputs(2170) <= (layer0_outputs(8474)) and not (layer0_outputs(6607));
    layer1_outputs(2171) <= (layer0_outputs(8920)) and not (layer0_outputs(8680));
    layer1_outputs(2172) <= not(layer0_outputs(7865)) or (layer0_outputs(6607));
    layer1_outputs(2173) <= not(layer0_outputs(422));
    layer1_outputs(2174) <= (layer0_outputs(3390)) xor (layer0_outputs(5990));
    layer1_outputs(2175) <= not((layer0_outputs(7258)) or (layer0_outputs(4657)));
    layer1_outputs(2176) <= layer0_outputs(8775);
    layer1_outputs(2177) <= '0';
    layer1_outputs(2178) <= not(layer0_outputs(6846));
    layer1_outputs(2179) <= (layer0_outputs(2450)) or (layer0_outputs(3264));
    layer1_outputs(2180) <= not((layer0_outputs(3958)) and (layer0_outputs(4045)));
    layer1_outputs(2181) <= (layer0_outputs(4030)) and (layer0_outputs(9835));
    layer1_outputs(2182) <= not(layer0_outputs(8430));
    layer1_outputs(2183) <= layer0_outputs(5418);
    layer1_outputs(2184) <= (layer0_outputs(6419)) and not (layer0_outputs(9023));
    layer1_outputs(2185) <= not(layer0_outputs(6284)) or (layer0_outputs(3634));
    layer1_outputs(2186) <= not(layer0_outputs(2677));
    layer1_outputs(2187) <= not(layer0_outputs(2292));
    layer1_outputs(2188) <= not((layer0_outputs(6771)) xor (layer0_outputs(6951)));
    layer1_outputs(2189) <= '0';
    layer1_outputs(2190) <= (layer0_outputs(9561)) and not (layer0_outputs(4649));
    layer1_outputs(2191) <= layer0_outputs(6727);
    layer1_outputs(2192) <= not((layer0_outputs(3515)) xor (layer0_outputs(1063)));
    layer1_outputs(2193) <= layer0_outputs(5738);
    layer1_outputs(2194) <= (layer0_outputs(5381)) and (layer0_outputs(2557));
    layer1_outputs(2195) <= not(layer0_outputs(8888));
    layer1_outputs(2196) <= not(layer0_outputs(6092));
    layer1_outputs(2197) <= layer0_outputs(10057);
    layer1_outputs(2198) <= (layer0_outputs(3116)) and not (layer0_outputs(6391));
    layer1_outputs(2199) <= (layer0_outputs(10202)) and (layer0_outputs(50));
    layer1_outputs(2200) <= not(layer0_outputs(1010));
    layer1_outputs(2201) <= not(layer0_outputs(7201)) or (layer0_outputs(5582));
    layer1_outputs(2202) <= (layer0_outputs(8801)) xor (layer0_outputs(3461));
    layer1_outputs(2203) <= not(layer0_outputs(6303));
    layer1_outputs(2204) <= layer0_outputs(8012);
    layer1_outputs(2205) <= not(layer0_outputs(311));
    layer1_outputs(2206) <= layer0_outputs(2303);
    layer1_outputs(2207) <= not(layer0_outputs(4022));
    layer1_outputs(2208) <= not(layer0_outputs(2013));
    layer1_outputs(2209) <= not(layer0_outputs(6042)) or (layer0_outputs(2291));
    layer1_outputs(2210) <= not(layer0_outputs(41));
    layer1_outputs(2211) <= not(layer0_outputs(9022));
    layer1_outputs(2212) <= not(layer0_outputs(5703));
    layer1_outputs(2213) <= not((layer0_outputs(1347)) or (layer0_outputs(4679)));
    layer1_outputs(2214) <= (layer0_outputs(8279)) and (layer0_outputs(6274));
    layer1_outputs(2215) <= (layer0_outputs(9013)) xor (layer0_outputs(770));
    layer1_outputs(2216) <= not((layer0_outputs(7485)) and (layer0_outputs(4)));
    layer1_outputs(2217) <= not((layer0_outputs(5219)) or (layer0_outputs(675)));
    layer1_outputs(2218) <= (layer0_outputs(9567)) or (layer0_outputs(1133));
    layer1_outputs(2219) <= '0';
    layer1_outputs(2220) <= (layer0_outputs(3912)) and not (layer0_outputs(6053));
    layer1_outputs(2221) <= not(layer0_outputs(8159));
    layer1_outputs(2222) <= not(layer0_outputs(6663));
    layer1_outputs(2223) <= layer0_outputs(590);
    layer1_outputs(2224) <= layer0_outputs(8981);
    layer1_outputs(2225) <= not(layer0_outputs(5425));
    layer1_outputs(2226) <= not(layer0_outputs(8251));
    layer1_outputs(2227) <= layer0_outputs(9267);
    layer1_outputs(2228) <= not(layer0_outputs(8528)) or (layer0_outputs(9758));
    layer1_outputs(2229) <= layer0_outputs(9554);
    layer1_outputs(2230) <= not((layer0_outputs(276)) and (layer0_outputs(3674)));
    layer1_outputs(2231) <= '1';
    layer1_outputs(2232) <= (layer0_outputs(2414)) and not (layer0_outputs(611));
    layer1_outputs(2233) <= not(layer0_outputs(1815)) or (layer0_outputs(570));
    layer1_outputs(2234) <= layer0_outputs(6127);
    layer1_outputs(2235) <= not(layer0_outputs(2315)) or (layer0_outputs(2761));
    layer1_outputs(2236) <= (layer0_outputs(4482)) and not (layer0_outputs(7762));
    layer1_outputs(2237) <= not(layer0_outputs(1053)) or (layer0_outputs(9311));
    layer1_outputs(2238) <= layer0_outputs(8176);
    layer1_outputs(2239) <= (layer0_outputs(4505)) and (layer0_outputs(5501));
    layer1_outputs(2240) <= (layer0_outputs(7909)) or (layer0_outputs(5052));
    layer1_outputs(2241) <= (layer0_outputs(104)) and not (layer0_outputs(683));
    layer1_outputs(2242) <= not(layer0_outputs(7108)) or (layer0_outputs(6318));
    layer1_outputs(2243) <= layer0_outputs(5958);
    layer1_outputs(2244) <= (layer0_outputs(4375)) and not (layer0_outputs(4337));
    layer1_outputs(2245) <= not(layer0_outputs(7717));
    layer1_outputs(2246) <= layer0_outputs(600);
    layer1_outputs(2247) <= not((layer0_outputs(8292)) or (layer0_outputs(6782)));
    layer1_outputs(2248) <= (layer0_outputs(3629)) and not (layer0_outputs(67));
    layer1_outputs(2249) <= not((layer0_outputs(432)) or (layer0_outputs(4435)));
    layer1_outputs(2250) <= (layer0_outputs(9602)) and not (layer0_outputs(8271));
    layer1_outputs(2251) <= (layer0_outputs(3542)) and not (layer0_outputs(1431));
    layer1_outputs(2252) <= (layer0_outputs(5938)) and not (layer0_outputs(6606));
    layer1_outputs(2253) <= (layer0_outputs(4218)) and (layer0_outputs(4624));
    layer1_outputs(2254) <= not(layer0_outputs(9527));
    layer1_outputs(2255) <= not((layer0_outputs(7340)) or (layer0_outputs(1083)));
    layer1_outputs(2256) <= not(layer0_outputs(8219));
    layer1_outputs(2257) <= not((layer0_outputs(5545)) xor (layer0_outputs(4411)));
    layer1_outputs(2258) <= layer0_outputs(5840);
    layer1_outputs(2259) <= not(layer0_outputs(3015));
    layer1_outputs(2260) <= (layer0_outputs(4222)) xor (layer0_outputs(8219));
    layer1_outputs(2261) <= not(layer0_outputs(6142)) or (layer0_outputs(2214));
    layer1_outputs(2262) <= (layer0_outputs(4162)) and not (layer0_outputs(48));
    layer1_outputs(2263) <= layer0_outputs(9633);
    layer1_outputs(2264) <= (layer0_outputs(6962)) and (layer0_outputs(4133));
    layer1_outputs(2265) <= not(layer0_outputs(2560));
    layer1_outputs(2266) <= layer0_outputs(8056);
    layer1_outputs(2267) <= not(layer0_outputs(9019));
    layer1_outputs(2268) <= not(layer0_outputs(5680)) or (layer0_outputs(9442));
    layer1_outputs(2269) <= layer0_outputs(6582);
    layer1_outputs(2270) <= not(layer0_outputs(60)) or (layer0_outputs(7397));
    layer1_outputs(2271) <= not(layer0_outputs(8194));
    layer1_outputs(2272) <= (layer0_outputs(3813)) xor (layer0_outputs(6745));
    layer1_outputs(2273) <= (layer0_outputs(9756)) xor (layer0_outputs(6253));
    layer1_outputs(2274) <= not(layer0_outputs(7730)) or (layer0_outputs(6074));
    layer1_outputs(2275) <= not((layer0_outputs(682)) and (layer0_outputs(1883)));
    layer1_outputs(2276) <= (layer0_outputs(425)) xor (layer0_outputs(5112));
    layer1_outputs(2277) <= (layer0_outputs(8975)) and not (layer0_outputs(7817));
    layer1_outputs(2278) <= layer0_outputs(974);
    layer1_outputs(2279) <= not(layer0_outputs(6928));
    layer1_outputs(2280) <= not((layer0_outputs(5944)) xor (layer0_outputs(4980)));
    layer1_outputs(2281) <= not(layer0_outputs(842)) or (layer0_outputs(56));
    layer1_outputs(2282) <= not(layer0_outputs(8374));
    layer1_outputs(2283) <= not(layer0_outputs(6815));
    layer1_outputs(2284) <= (layer0_outputs(1037)) xor (layer0_outputs(4470));
    layer1_outputs(2285) <= layer0_outputs(6372);
    layer1_outputs(2286) <= (layer0_outputs(7203)) or (layer0_outputs(8445));
    layer1_outputs(2287) <= layer0_outputs(7897);
    layer1_outputs(2288) <= not(layer0_outputs(8001)) or (layer0_outputs(6142));
    layer1_outputs(2289) <= not((layer0_outputs(5333)) or (layer0_outputs(576)));
    layer1_outputs(2290) <= (layer0_outputs(6703)) xor (layer0_outputs(2164));
    layer1_outputs(2291) <= (layer0_outputs(3779)) and (layer0_outputs(837));
    layer1_outputs(2292) <= layer0_outputs(4172);
    layer1_outputs(2293) <= (layer0_outputs(9101)) and not (layer0_outputs(8156));
    layer1_outputs(2294) <= not(layer0_outputs(4799));
    layer1_outputs(2295) <= not(layer0_outputs(5636));
    layer1_outputs(2296) <= not(layer0_outputs(4624)) or (layer0_outputs(90));
    layer1_outputs(2297) <= not(layer0_outputs(2126)) or (layer0_outputs(3169));
    layer1_outputs(2298) <= (layer0_outputs(7191)) or (layer0_outputs(6220));
    layer1_outputs(2299) <= not(layer0_outputs(9834)) or (layer0_outputs(8193));
    layer1_outputs(2300) <= not((layer0_outputs(9173)) or (layer0_outputs(5760)));
    layer1_outputs(2301) <= (layer0_outputs(7258)) and not (layer0_outputs(8115));
    layer1_outputs(2302) <= layer0_outputs(6216);
    layer1_outputs(2303) <= not(layer0_outputs(4104));
    layer1_outputs(2304) <= not(layer0_outputs(4138));
    layer1_outputs(2305) <= not((layer0_outputs(9841)) and (layer0_outputs(239)));
    layer1_outputs(2306) <= not((layer0_outputs(942)) xor (layer0_outputs(1595)));
    layer1_outputs(2307) <= not((layer0_outputs(4623)) xor (layer0_outputs(3503)));
    layer1_outputs(2308) <= (layer0_outputs(7005)) and not (layer0_outputs(3429));
    layer1_outputs(2309) <= not((layer0_outputs(5001)) and (layer0_outputs(8683)));
    layer1_outputs(2310) <= not(layer0_outputs(8590)) or (layer0_outputs(4121));
    layer1_outputs(2311) <= (layer0_outputs(7708)) xor (layer0_outputs(9480));
    layer1_outputs(2312) <= not(layer0_outputs(5810));
    layer1_outputs(2313) <= (layer0_outputs(1935)) or (layer0_outputs(691));
    layer1_outputs(2314) <= not((layer0_outputs(5398)) and (layer0_outputs(2566)));
    layer1_outputs(2315) <= not(layer0_outputs(5665)) or (layer0_outputs(5256));
    layer1_outputs(2316) <= not((layer0_outputs(6316)) or (layer0_outputs(2471)));
    layer1_outputs(2317) <= not((layer0_outputs(7221)) and (layer0_outputs(6031)));
    layer1_outputs(2318) <= not((layer0_outputs(9496)) and (layer0_outputs(1044)));
    layer1_outputs(2319) <= (layer0_outputs(3891)) and not (layer0_outputs(7152));
    layer1_outputs(2320) <= (layer0_outputs(3186)) and not (layer0_outputs(3503));
    layer1_outputs(2321) <= not((layer0_outputs(4296)) xor (layer0_outputs(4591)));
    layer1_outputs(2322) <= (layer0_outputs(5735)) or (layer0_outputs(3687));
    layer1_outputs(2323) <= layer0_outputs(10008);
    layer1_outputs(2324) <= (layer0_outputs(1716)) and not (layer0_outputs(9062));
    layer1_outputs(2325) <= not(layer0_outputs(3221));
    layer1_outputs(2326) <= not((layer0_outputs(5)) xor (layer0_outputs(7725)));
    layer1_outputs(2327) <= not((layer0_outputs(2807)) or (layer0_outputs(2975)));
    layer1_outputs(2328) <= not(layer0_outputs(7066)) or (layer0_outputs(8707));
    layer1_outputs(2329) <= not(layer0_outputs(8003)) or (layer0_outputs(861));
    layer1_outputs(2330) <= layer0_outputs(2710);
    layer1_outputs(2331) <= (layer0_outputs(591)) and not (layer0_outputs(7874));
    layer1_outputs(2332) <= layer0_outputs(9971);
    layer1_outputs(2333) <= not(layer0_outputs(6978));
    layer1_outputs(2334) <= not(layer0_outputs(9803)) or (layer0_outputs(7999));
    layer1_outputs(2335) <= not(layer0_outputs(6768));
    layer1_outputs(2336) <= '1';
    layer1_outputs(2337) <= layer0_outputs(2169);
    layer1_outputs(2338) <= not((layer0_outputs(5138)) xor (layer0_outputs(7972)));
    layer1_outputs(2339) <= (layer0_outputs(2936)) xor (layer0_outputs(5705));
    layer1_outputs(2340) <= not((layer0_outputs(7442)) and (layer0_outputs(4688)));
    layer1_outputs(2341) <= (layer0_outputs(9589)) and (layer0_outputs(1970));
    layer1_outputs(2342) <= not(layer0_outputs(6559));
    layer1_outputs(2343) <= not(layer0_outputs(2101));
    layer1_outputs(2344) <= layer0_outputs(642);
    layer1_outputs(2345) <= layer0_outputs(2966);
    layer1_outputs(2346) <= layer0_outputs(8925);
    layer1_outputs(2347) <= layer0_outputs(549);
    layer1_outputs(2348) <= not((layer0_outputs(253)) and (layer0_outputs(546)));
    layer1_outputs(2349) <= layer0_outputs(9558);
    layer1_outputs(2350) <= layer0_outputs(8979);
    layer1_outputs(2351) <= not(layer0_outputs(626));
    layer1_outputs(2352) <= '0';
    layer1_outputs(2353) <= not(layer0_outputs(3081)) or (layer0_outputs(2098));
    layer1_outputs(2354) <= not(layer0_outputs(4052)) or (layer0_outputs(1038));
    layer1_outputs(2355) <= not((layer0_outputs(9379)) or (layer0_outputs(5480)));
    layer1_outputs(2356) <= layer0_outputs(5767);
    layer1_outputs(2357) <= layer0_outputs(9870);
    layer1_outputs(2358) <= (layer0_outputs(7334)) and not (layer0_outputs(3329));
    layer1_outputs(2359) <= not((layer0_outputs(7756)) or (layer0_outputs(4089)));
    layer1_outputs(2360) <= not((layer0_outputs(9597)) and (layer0_outputs(1951)));
    layer1_outputs(2361) <= not((layer0_outputs(2615)) xor (layer0_outputs(6344)));
    layer1_outputs(2362) <= not(layer0_outputs(4677));
    layer1_outputs(2363) <= not(layer0_outputs(3146)) or (layer0_outputs(3635));
    layer1_outputs(2364) <= not(layer0_outputs(9564));
    layer1_outputs(2365) <= layer0_outputs(6181);
    layer1_outputs(2366) <= (layer0_outputs(4907)) and (layer0_outputs(5376));
    layer1_outputs(2367) <= not(layer0_outputs(508));
    layer1_outputs(2368) <= layer0_outputs(3297);
    layer1_outputs(2369) <= not(layer0_outputs(6156));
    layer1_outputs(2370) <= not(layer0_outputs(9385)) or (layer0_outputs(2974));
    layer1_outputs(2371) <= not(layer0_outputs(4724)) or (layer0_outputs(7806));
    layer1_outputs(2372) <= not((layer0_outputs(1479)) and (layer0_outputs(6276)));
    layer1_outputs(2373) <= not(layer0_outputs(8062));
    layer1_outputs(2374) <= not((layer0_outputs(8853)) or (layer0_outputs(2599)));
    layer1_outputs(2375) <= (layer0_outputs(5210)) and not (layer0_outputs(2544));
    layer1_outputs(2376) <= not(layer0_outputs(3153));
    layer1_outputs(2377) <= (layer0_outputs(2657)) and not (layer0_outputs(6941));
    layer1_outputs(2378) <= '1';
    layer1_outputs(2379) <= (layer0_outputs(1093)) and not (layer0_outputs(6306));
    layer1_outputs(2380) <= not(layer0_outputs(3331));
    layer1_outputs(2381) <= layer0_outputs(4082);
    layer1_outputs(2382) <= (layer0_outputs(1458)) xor (layer0_outputs(4020));
    layer1_outputs(2383) <= not(layer0_outputs(2118)) or (layer0_outputs(4966));
    layer1_outputs(2384) <= not(layer0_outputs(1343));
    layer1_outputs(2385) <= not((layer0_outputs(1269)) xor (layer0_outputs(8660)));
    layer1_outputs(2386) <= (layer0_outputs(9735)) or (layer0_outputs(3137));
    layer1_outputs(2387) <= not((layer0_outputs(9211)) and (layer0_outputs(6944)));
    layer1_outputs(2388) <= (layer0_outputs(7138)) and (layer0_outputs(9057));
    layer1_outputs(2389) <= not((layer0_outputs(7095)) xor (layer0_outputs(5825)));
    layer1_outputs(2390) <= not(layer0_outputs(4381));
    layer1_outputs(2391) <= not(layer0_outputs(7310)) or (layer0_outputs(5963));
    layer1_outputs(2392) <= layer0_outputs(3420);
    layer1_outputs(2393) <= not((layer0_outputs(6505)) xor (layer0_outputs(8767)));
    layer1_outputs(2394) <= not(layer0_outputs(7751)) or (layer0_outputs(3538));
    layer1_outputs(2395) <= '1';
    layer1_outputs(2396) <= not(layer0_outputs(7316)) or (layer0_outputs(5569));
    layer1_outputs(2397) <= not((layer0_outputs(2307)) xor (layer0_outputs(314)));
    layer1_outputs(2398) <= not((layer0_outputs(8002)) and (layer0_outputs(6390)));
    layer1_outputs(2399) <= layer0_outputs(7854);
    layer1_outputs(2400) <= not(layer0_outputs(9880));
    layer1_outputs(2401) <= not((layer0_outputs(4511)) and (layer0_outputs(5039)));
    layer1_outputs(2402) <= not(layer0_outputs(3444)) or (layer0_outputs(8535));
    layer1_outputs(2403) <= '0';
    layer1_outputs(2404) <= (layer0_outputs(2711)) xor (layer0_outputs(4582));
    layer1_outputs(2405) <= (layer0_outputs(9443)) and not (layer0_outputs(3198));
    layer1_outputs(2406) <= not(layer0_outputs(7271));
    layer1_outputs(2407) <= layer0_outputs(3560);
    layer1_outputs(2408) <= (layer0_outputs(6629)) xor (layer0_outputs(3487));
    layer1_outputs(2409) <= (layer0_outputs(4832)) and (layer0_outputs(6603));
    layer1_outputs(2410) <= not(layer0_outputs(666)) or (layer0_outputs(8616));
    layer1_outputs(2411) <= not(layer0_outputs(3195));
    layer1_outputs(2412) <= layer0_outputs(642);
    layer1_outputs(2413) <= not((layer0_outputs(2692)) or (layer0_outputs(7215)));
    layer1_outputs(2414) <= (layer0_outputs(354)) xor (layer0_outputs(9217));
    layer1_outputs(2415) <= (layer0_outputs(9592)) or (layer0_outputs(6175));
    layer1_outputs(2416) <= not((layer0_outputs(7884)) and (layer0_outputs(5137)));
    layer1_outputs(2417) <= (layer0_outputs(9193)) and not (layer0_outputs(5441));
    layer1_outputs(2418) <= (layer0_outputs(505)) xor (layer0_outputs(5015));
    layer1_outputs(2419) <= not(layer0_outputs(868));
    layer1_outputs(2420) <= (layer0_outputs(8226)) and (layer0_outputs(9534));
    layer1_outputs(2421) <= not((layer0_outputs(3596)) and (layer0_outputs(5001)));
    layer1_outputs(2422) <= (layer0_outputs(9143)) and not (layer0_outputs(4369));
    layer1_outputs(2423) <= not(layer0_outputs(9489)) or (layer0_outputs(2855));
    layer1_outputs(2424) <= layer0_outputs(7584);
    layer1_outputs(2425) <= layer0_outputs(723);
    layer1_outputs(2426) <= (layer0_outputs(6751)) and (layer0_outputs(9812));
    layer1_outputs(2427) <= (layer0_outputs(944)) xor (layer0_outputs(1640));
    layer1_outputs(2428) <= not((layer0_outputs(5318)) and (layer0_outputs(3042)));
    layer1_outputs(2429) <= not(layer0_outputs(3205));
    layer1_outputs(2430) <= not(layer0_outputs(1941)) or (layer0_outputs(9950));
    layer1_outputs(2431) <= not((layer0_outputs(2655)) or (layer0_outputs(847)));
    layer1_outputs(2432) <= (layer0_outputs(7506)) xor (layer0_outputs(3109));
    layer1_outputs(2433) <= (layer0_outputs(2817)) or (layer0_outputs(6018));
    layer1_outputs(2434) <= layer0_outputs(8339);
    layer1_outputs(2435) <= not(layer0_outputs(2852));
    layer1_outputs(2436) <= layer0_outputs(6255);
    layer1_outputs(2437) <= (layer0_outputs(5204)) and (layer0_outputs(4436));
    layer1_outputs(2438) <= '1';
    layer1_outputs(2439) <= layer0_outputs(5481);
    layer1_outputs(2440) <= (layer0_outputs(141)) or (layer0_outputs(10041));
    layer1_outputs(2441) <= (layer0_outputs(9818)) and (layer0_outputs(7270));
    layer1_outputs(2442) <= not((layer0_outputs(1818)) and (layer0_outputs(1104)));
    layer1_outputs(2443) <= not(layer0_outputs(8898));
    layer1_outputs(2444) <= (layer0_outputs(3941)) and not (layer0_outputs(3277));
    layer1_outputs(2445) <= layer0_outputs(9737);
    layer1_outputs(2446) <= (layer0_outputs(8940)) xor (layer0_outputs(5293));
    layer1_outputs(2447) <= (layer0_outputs(6937)) xor (layer0_outputs(6500));
    layer1_outputs(2448) <= '1';
    layer1_outputs(2449) <= layer0_outputs(1446);
    layer1_outputs(2450) <= layer0_outputs(2534);
    layer1_outputs(2451) <= not((layer0_outputs(2981)) or (layer0_outputs(1275)));
    layer1_outputs(2452) <= layer0_outputs(6962);
    layer1_outputs(2453) <= layer0_outputs(5608);
    layer1_outputs(2454) <= not((layer0_outputs(9501)) and (layer0_outputs(3184)));
    layer1_outputs(2455) <= layer0_outputs(8074);
    layer1_outputs(2456) <= '1';
    layer1_outputs(2457) <= not((layer0_outputs(6704)) or (layer0_outputs(9072)));
    layer1_outputs(2458) <= not(layer0_outputs(9595));
    layer1_outputs(2459) <= (layer0_outputs(8095)) and (layer0_outputs(9796));
    layer1_outputs(2460) <= (layer0_outputs(8666)) and not (layer0_outputs(7249));
    layer1_outputs(2461) <= not(layer0_outputs(7227)) or (layer0_outputs(1516));
    layer1_outputs(2462) <= (layer0_outputs(4146)) xor (layer0_outputs(8756));
    layer1_outputs(2463) <= (layer0_outputs(1700)) or (layer0_outputs(9360));
    layer1_outputs(2464) <= layer0_outputs(5775);
    layer1_outputs(2465) <= (layer0_outputs(9901)) or (layer0_outputs(9158));
    layer1_outputs(2466) <= not(layer0_outputs(1061)) or (layer0_outputs(7314));
    layer1_outputs(2467) <= layer0_outputs(2176);
    layer1_outputs(2468) <= (layer0_outputs(7550)) and not (layer0_outputs(9268));
    layer1_outputs(2469) <= layer0_outputs(7869);
    layer1_outputs(2470) <= not(layer0_outputs(8682));
    layer1_outputs(2471) <= not((layer0_outputs(4146)) or (layer0_outputs(8055)));
    layer1_outputs(2472) <= not((layer0_outputs(8674)) and (layer0_outputs(3299)));
    layer1_outputs(2473) <= layer0_outputs(4737);
    layer1_outputs(2474) <= (layer0_outputs(7709)) xor (layer0_outputs(9506));
    layer1_outputs(2475) <= (layer0_outputs(152)) xor (layer0_outputs(8476));
    layer1_outputs(2476) <= not(layer0_outputs(7441)) or (layer0_outputs(1366));
    layer1_outputs(2477) <= not(layer0_outputs(8667));
    layer1_outputs(2478) <= layer0_outputs(6983);
    layer1_outputs(2479) <= (layer0_outputs(8759)) and not (layer0_outputs(4784));
    layer1_outputs(2480) <= not((layer0_outputs(4134)) and (layer0_outputs(4409)));
    layer1_outputs(2481) <= layer0_outputs(8752);
    layer1_outputs(2482) <= not(layer0_outputs(808));
    layer1_outputs(2483) <= (layer0_outputs(2434)) and not (layer0_outputs(6223));
    layer1_outputs(2484) <= not(layer0_outputs(8149));
    layer1_outputs(2485) <= not((layer0_outputs(1534)) xor (layer0_outputs(7118)));
    layer1_outputs(2486) <= (layer0_outputs(9548)) and not (layer0_outputs(5092));
    layer1_outputs(2487) <= not(layer0_outputs(6555));
    layer1_outputs(2488) <= layer0_outputs(2297);
    layer1_outputs(2489) <= not((layer0_outputs(8048)) or (layer0_outputs(9276)));
    layer1_outputs(2490) <= not(layer0_outputs(5817));
    layer1_outputs(2491) <= not((layer0_outputs(8333)) or (layer0_outputs(230)));
    layer1_outputs(2492) <= (layer0_outputs(10186)) or (layer0_outputs(8105));
    layer1_outputs(2493) <= (layer0_outputs(1440)) and not (layer0_outputs(6546));
    layer1_outputs(2494) <= layer0_outputs(6458);
    layer1_outputs(2495) <= (layer0_outputs(9053)) and (layer0_outputs(6953));
    layer1_outputs(2496) <= (layer0_outputs(3821)) and not (layer0_outputs(1514));
    layer1_outputs(2497) <= layer0_outputs(4165);
    layer1_outputs(2498) <= (layer0_outputs(7345)) and (layer0_outputs(2666));
    layer1_outputs(2499) <= not((layer0_outputs(3874)) xor (layer0_outputs(8419)));
    layer1_outputs(2500) <= layer0_outputs(8249);
    layer1_outputs(2501) <= not(layer0_outputs(3630)) or (layer0_outputs(8956));
    layer1_outputs(2502) <= not(layer0_outputs(3291));
    layer1_outputs(2503) <= layer0_outputs(5819);
    layer1_outputs(2504) <= not(layer0_outputs(7889)) or (layer0_outputs(5043));
    layer1_outputs(2505) <= layer0_outputs(1878);
    layer1_outputs(2506) <= not((layer0_outputs(8183)) or (layer0_outputs(7345)));
    layer1_outputs(2507) <= not((layer0_outputs(9165)) and (layer0_outputs(5741)));
    layer1_outputs(2508) <= layer0_outputs(5260);
    layer1_outputs(2509) <= (layer0_outputs(3180)) and not (layer0_outputs(4415));
    layer1_outputs(2510) <= layer0_outputs(1307);
    layer1_outputs(2511) <= not(layer0_outputs(6707)) or (layer0_outputs(3296));
    layer1_outputs(2512) <= layer0_outputs(10179);
    layer1_outputs(2513) <= layer0_outputs(5251);
    layer1_outputs(2514) <= layer0_outputs(9850);
    layer1_outputs(2515) <= (layer0_outputs(7619)) xor (layer0_outputs(9640));
    layer1_outputs(2516) <= not(layer0_outputs(5771));
    layer1_outputs(2517) <= not(layer0_outputs(2162)) or (layer0_outputs(42));
    layer1_outputs(2518) <= layer0_outputs(10080);
    layer1_outputs(2519) <= not(layer0_outputs(2847));
    layer1_outputs(2520) <= layer0_outputs(7197);
    layer1_outputs(2521) <= (layer0_outputs(6702)) xor (layer0_outputs(1214));
    layer1_outputs(2522) <= not(layer0_outputs(9382)) or (layer0_outputs(8310));
    layer1_outputs(2523) <= layer0_outputs(9690);
    layer1_outputs(2524) <= not((layer0_outputs(1071)) and (layer0_outputs(5163)));
    layer1_outputs(2525) <= not(layer0_outputs(1740)) or (layer0_outputs(1685));
    layer1_outputs(2526) <= (layer0_outputs(5489)) and not (layer0_outputs(7702));
    layer1_outputs(2527) <= (layer0_outputs(542)) and (layer0_outputs(3352));
    layer1_outputs(2528) <= not(layer0_outputs(6839));
    layer1_outputs(2529) <= (layer0_outputs(8626)) and (layer0_outputs(414));
    layer1_outputs(2530) <= (layer0_outputs(3726)) and not (layer0_outputs(3474));
    layer1_outputs(2531) <= (layer0_outputs(703)) xor (layer0_outputs(1521));
    layer1_outputs(2532) <= not(layer0_outputs(4073)) or (layer0_outputs(5102));
    layer1_outputs(2533) <= layer0_outputs(797);
    layer1_outputs(2534) <= not(layer0_outputs(8338));
    layer1_outputs(2535) <= not((layer0_outputs(687)) xor (layer0_outputs(2255)));
    layer1_outputs(2536) <= layer0_outputs(3395);
    layer1_outputs(2537) <= not(layer0_outputs(8564));
    layer1_outputs(2538) <= (layer0_outputs(6450)) or (layer0_outputs(3203));
    layer1_outputs(2539) <= (layer0_outputs(7128)) xor (layer0_outputs(3119));
    layer1_outputs(2540) <= layer0_outputs(7214);
    layer1_outputs(2541) <= layer0_outputs(8055);
    layer1_outputs(2542) <= not((layer0_outputs(9905)) and (layer0_outputs(3100)));
    layer1_outputs(2543) <= layer0_outputs(1306);
    layer1_outputs(2544) <= layer0_outputs(2987);
    layer1_outputs(2545) <= layer0_outputs(654);
    layer1_outputs(2546) <= not(layer0_outputs(3606));
    layer1_outputs(2547) <= not(layer0_outputs(74)) or (layer0_outputs(8417));
    layer1_outputs(2548) <= layer0_outputs(3062);
    layer1_outputs(2549) <= not(layer0_outputs(9343));
    layer1_outputs(2550) <= not(layer0_outputs(6904)) or (layer0_outputs(2983));
    layer1_outputs(2551) <= (layer0_outputs(9433)) or (layer0_outputs(7474));
    layer1_outputs(2552) <= layer0_outputs(4332);
    layer1_outputs(2553) <= layer0_outputs(8530);
    layer1_outputs(2554) <= (layer0_outputs(7558)) xor (layer0_outputs(5534));
    layer1_outputs(2555) <= (layer0_outputs(6307)) and (layer0_outputs(2524));
    layer1_outputs(2556) <= not(layer0_outputs(9719));
    layer1_outputs(2557) <= layer0_outputs(5962);
    layer1_outputs(2558) <= not(layer0_outputs(9463)) or (layer0_outputs(376));
    layer1_outputs(2559) <= (layer0_outputs(5596)) and not (layer0_outputs(4956));
    layer1_outputs(2560) <= not((layer0_outputs(51)) and (layer0_outputs(6105)));
    layer1_outputs(2561) <= layer0_outputs(7387);
    layer1_outputs(2562) <= (layer0_outputs(9621)) and not (layer0_outputs(9837));
    layer1_outputs(2563) <= layer0_outputs(5207);
    layer1_outputs(2564) <= layer0_outputs(4764);
    layer1_outputs(2565) <= not((layer0_outputs(1432)) or (layer0_outputs(9977)));
    layer1_outputs(2566) <= (layer0_outputs(1362)) and not (layer0_outputs(4562));
    layer1_outputs(2567) <= (layer0_outputs(8554)) or (layer0_outputs(7024));
    layer1_outputs(2568) <= not(layer0_outputs(5661));
    layer1_outputs(2569) <= not(layer0_outputs(10094));
    layer1_outputs(2570) <= (layer0_outputs(1254)) and not (layer0_outputs(7507));
    layer1_outputs(2571) <= (layer0_outputs(7698)) and not (layer0_outputs(9780));
    layer1_outputs(2572) <= not(layer0_outputs(2106));
    layer1_outputs(2573) <= not(layer0_outputs(745)) or (layer0_outputs(2740));
    layer1_outputs(2574) <= layer0_outputs(6046);
    layer1_outputs(2575) <= (layer0_outputs(5028)) and not (layer0_outputs(5448));
    layer1_outputs(2576) <= not(layer0_outputs(7594)) or (layer0_outputs(2253));
    layer1_outputs(2577) <= (layer0_outputs(1320)) and (layer0_outputs(8806));
    layer1_outputs(2578) <= (layer0_outputs(3215)) xor (layer0_outputs(3522));
    layer1_outputs(2579) <= not((layer0_outputs(7124)) or (layer0_outputs(9857)));
    layer1_outputs(2580) <= layer0_outputs(4919);
    layer1_outputs(2581) <= not((layer0_outputs(1449)) and (layer0_outputs(8093)));
    layer1_outputs(2582) <= not(layer0_outputs(1478)) or (layer0_outputs(3727));
    layer1_outputs(2583) <= not(layer0_outputs(945));
    layer1_outputs(2584) <= not(layer0_outputs(4293));
    layer1_outputs(2585) <= not((layer0_outputs(6795)) xor (layer0_outputs(2087)));
    layer1_outputs(2586) <= '0';
    layer1_outputs(2587) <= not(layer0_outputs(9111));
    layer1_outputs(2588) <= not(layer0_outputs(462));
    layer1_outputs(2589) <= not(layer0_outputs(1092)) or (layer0_outputs(9896));
    layer1_outputs(2590) <= not(layer0_outputs(2716));
    layer1_outputs(2591) <= (layer0_outputs(7575)) and (layer0_outputs(8737));
    layer1_outputs(2592) <= not(layer0_outputs(9249));
    layer1_outputs(2593) <= not((layer0_outputs(8379)) and (layer0_outputs(8122)));
    layer1_outputs(2594) <= not(layer0_outputs(887)) or (layer0_outputs(1930));
    layer1_outputs(2595) <= not(layer0_outputs(993));
    layer1_outputs(2596) <= layer0_outputs(9752);
    layer1_outputs(2597) <= not((layer0_outputs(310)) and (layer0_outputs(1478)));
    layer1_outputs(2598) <= layer0_outputs(10197);
    layer1_outputs(2599) <= layer0_outputs(5654);
    layer1_outputs(2600) <= not((layer0_outputs(9593)) xor (layer0_outputs(3359)));
    layer1_outputs(2601) <= layer0_outputs(4857);
    layer1_outputs(2602) <= not(layer0_outputs(3265));
    layer1_outputs(2603) <= not((layer0_outputs(1032)) xor (layer0_outputs(5181)));
    layer1_outputs(2604) <= not((layer0_outputs(4918)) xor (layer0_outputs(2312)));
    layer1_outputs(2605) <= not((layer0_outputs(1278)) xor (layer0_outputs(3424)));
    layer1_outputs(2606) <= not((layer0_outputs(6218)) xor (layer0_outputs(5896)));
    layer1_outputs(2607) <= not((layer0_outputs(10094)) or (layer0_outputs(4571)));
    layer1_outputs(2608) <= not(layer0_outputs(7261)) or (layer0_outputs(8915));
    layer1_outputs(2609) <= layer0_outputs(1592);
    layer1_outputs(2610) <= not(layer0_outputs(6661)) or (layer0_outputs(2721));
    layer1_outputs(2611) <= not(layer0_outputs(6794));
    layer1_outputs(2612) <= not(layer0_outputs(1735));
    layer1_outputs(2613) <= not(layer0_outputs(3857));
    layer1_outputs(2614) <= not(layer0_outputs(9292));
    layer1_outputs(2615) <= (layer0_outputs(5621)) and not (layer0_outputs(5394));
    layer1_outputs(2616) <= layer0_outputs(841);
    layer1_outputs(2617) <= layer0_outputs(2202);
    layer1_outputs(2618) <= not(layer0_outputs(6695));
    layer1_outputs(2619) <= layer0_outputs(5118);
    layer1_outputs(2620) <= (layer0_outputs(5755)) xor (layer0_outputs(503));
    layer1_outputs(2621) <= (layer0_outputs(2487)) or (layer0_outputs(2065));
    layer1_outputs(2622) <= layer0_outputs(9518);
    layer1_outputs(2623) <= layer0_outputs(5232);
    layer1_outputs(2624) <= not((layer0_outputs(7802)) xor (layer0_outputs(9410)));
    layer1_outputs(2625) <= layer0_outputs(6928);
    layer1_outputs(2626) <= (layer0_outputs(871)) or (layer0_outputs(6088));
    layer1_outputs(2627) <= not((layer0_outputs(1099)) or (layer0_outputs(6331)));
    layer1_outputs(2628) <= '1';
    layer1_outputs(2629) <= not((layer0_outputs(8830)) or (layer0_outputs(2295)));
    layer1_outputs(2630) <= not(layer0_outputs(6240)) or (layer0_outputs(1434));
    layer1_outputs(2631) <= layer0_outputs(9307);
    layer1_outputs(2632) <= layer0_outputs(5558);
    layer1_outputs(2633) <= (layer0_outputs(8777)) and (layer0_outputs(5163));
    layer1_outputs(2634) <= layer0_outputs(1812);
    layer1_outputs(2635) <= not((layer0_outputs(8709)) xor (layer0_outputs(6461)));
    layer1_outputs(2636) <= (layer0_outputs(3054)) or (layer0_outputs(3505));
    layer1_outputs(2637) <= not((layer0_outputs(8239)) or (layer0_outputs(1013)));
    layer1_outputs(2638) <= layer0_outputs(9567);
    layer1_outputs(2639) <= not((layer0_outputs(4013)) or (layer0_outputs(6131)));
    layer1_outputs(2640) <= not(layer0_outputs(6999));
    layer1_outputs(2641) <= not((layer0_outputs(9267)) or (layer0_outputs(4748)));
    layer1_outputs(2642) <= layer0_outputs(2478);
    layer1_outputs(2643) <= layer0_outputs(5691);
    layer1_outputs(2644) <= (layer0_outputs(2117)) and not (layer0_outputs(2447));
    layer1_outputs(2645) <= '0';
    layer1_outputs(2646) <= '0';
    layer1_outputs(2647) <= not(layer0_outputs(9322)) or (layer0_outputs(5573));
    layer1_outputs(2648) <= not((layer0_outputs(8388)) or (layer0_outputs(2860)));
    layer1_outputs(2649) <= (layer0_outputs(6299)) xor (layer0_outputs(1544));
    layer1_outputs(2650) <= not((layer0_outputs(5054)) or (layer0_outputs(705)));
    layer1_outputs(2651) <= layer0_outputs(6767);
    layer1_outputs(2652) <= not(layer0_outputs(7236));
    layer1_outputs(2653) <= not(layer0_outputs(5525)) or (layer0_outputs(8134));
    layer1_outputs(2654) <= (layer0_outputs(9597)) and not (layer0_outputs(6497));
    layer1_outputs(2655) <= (layer0_outputs(8078)) and not (layer0_outputs(6298));
    layer1_outputs(2656) <= (layer0_outputs(6467)) and (layer0_outputs(6759));
    layer1_outputs(2657) <= layer0_outputs(5997);
    layer1_outputs(2658) <= (layer0_outputs(1578)) or (layer0_outputs(6612));
    layer1_outputs(2659) <= layer0_outputs(4790);
    layer1_outputs(2660) <= not(layer0_outputs(7115));
    layer1_outputs(2661) <= layer0_outputs(1778);
    layer1_outputs(2662) <= (layer0_outputs(3040)) or (layer0_outputs(7424));
    layer1_outputs(2663) <= not((layer0_outputs(2296)) and (layer0_outputs(6026)));
    layer1_outputs(2664) <= (layer0_outputs(6237)) and (layer0_outputs(6598));
    layer1_outputs(2665) <= not(layer0_outputs(7211));
    layer1_outputs(2666) <= (layer0_outputs(1515)) and not (layer0_outputs(3310));
    layer1_outputs(2667) <= not(layer0_outputs(5554)) or (layer0_outputs(5333));
    layer1_outputs(2668) <= (layer0_outputs(2224)) and (layer0_outputs(6754));
    layer1_outputs(2669) <= not((layer0_outputs(7129)) and (layer0_outputs(9794)));
    layer1_outputs(2670) <= not(layer0_outputs(8617));
    layer1_outputs(2671) <= not((layer0_outputs(2997)) and (layer0_outputs(5082)));
    layer1_outputs(2672) <= (layer0_outputs(560)) and not (layer0_outputs(1126));
    layer1_outputs(2673) <= layer0_outputs(8161);
    layer1_outputs(2674) <= not((layer0_outputs(4612)) and (layer0_outputs(4421)));
    layer1_outputs(2675) <= not(layer0_outputs(9706));
    layer1_outputs(2676) <= (layer0_outputs(6252)) and not (layer0_outputs(3729));
    layer1_outputs(2677) <= not(layer0_outputs(4714));
    layer1_outputs(2678) <= not((layer0_outputs(9906)) xor (layer0_outputs(3823)));
    layer1_outputs(2679) <= not(layer0_outputs(4059)) or (layer0_outputs(4468));
    layer1_outputs(2680) <= layer0_outputs(7176);
    layer1_outputs(2681) <= (layer0_outputs(3086)) or (layer0_outputs(3670));
    layer1_outputs(2682) <= layer0_outputs(7328);
    layer1_outputs(2683) <= layer0_outputs(4704);
    layer1_outputs(2684) <= not(layer0_outputs(656)) or (layer0_outputs(224));
    layer1_outputs(2685) <= not(layer0_outputs(6323)) or (layer0_outputs(940));
    layer1_outputs(2686) <= '1';
    layer1_outputs(2687) <= not(layer0_outputs(738)) or (layer0_outputs(2072));
    layer1_outputs(2688) <= not((layer0_outputs(7297)) and (layer0_outputs(3849)));
    layer1_outputs(2689) <= layer0_outputs(8865);
    layer1_outputs(2690) <= not(layer0_outputs(6521));
    layer1_outputs(2691) <= layer0_outputs(1274);
    layer1_outputs(2692) <= not((layer0_outputs(6586)) and (layer0_outputs(5450)));
    layer1_outputs(2693) <= not(layer0_outputs(7626)) or (layer0_outputs(8822));
    layer1_outputs(2694) <= (layer0_outputs(5831)) or (layer0_outputs(1135));
    layer1_outputs(2695) <= not(layer0_outputs(2096));
    layer1_outputs(2696) <= (layer0_outputs(869)) and not (layer0_outputs(2813));
    layer1_outputs(2697) <= (layer0_outputs(7228)) or (layer0_outputs(7313));
    layer1_outputs(2698) <= layer0_outputs(9664);
    layer1_outputs(2699) <= (layer0_outputs(133)) xor (layer0_outputs(5505));
    layer1_outputs(2700) <= layer0_outputs(4114);
    layer1_outputs(2701) <= layer0_outputs(5443);
    layer1_outputs(2702) <= not(layer0_outputs(3876));
    layer1_outputs(2703) <= not(layer0_outputs(841)) or (layer0_outputs(6722));
    layer1_outputs(2704) <= not(layer0_outputs(9397)) or (layer0_outputs(2366));
    layer1_outputs(2705) <= not(layer0_outputs(4640)) or (layer0_outputs(6557));
    layer1_outputs(2706) <= not((layer0_outputs(7446)) or (layer0_outputs(5299)));
    layer1_outputs(2707) <= layer0_outputs(5391);
    layer1_outputs(2708) <= not(layer0_outputs(1337));
    layer1_outputs(2709) <= not(layer0_outputs(934));
    layer1_outputs(2710) <= not(layer0_outputs(4215));
    layer1_outputs(2711) <= not((layer0_outputs(7231)) or (layer0_outputs(3381)));
    layer1_outputs(2712) <= (layer0_outputs(4165)) and (layer0_outputs(4898));
    layer1_outputs(2713) <= '1';
    layer1_outputs(2714) <= layer0_outputs(371);
    layer1_outputs(2715) <= not((layer0_outputs(5511)) and (layer0_outputs(2408)));
    layer1_outputs(2716) <= not((layer0_outputs(7373)) and (layer0_outputs(680)));
    layer1_outputs(2717) <= not(layer0_outputs(9222)) or (layer0_outputs(648));
    layer1_outputs(2718) <= not(layer0_outputs(4005)) or (layer0_outputs(2002));
    layer1_outputs(2719) <= not((layer0_outputs(4023)) xor (layer0_outputs(5404)));
    layer1_outputs(2720) <= '0';
    layer1_outputs(2721) <= layer0_outputs(5472);
    layer1_outputs(2722) <= not((layer0_outputs(3894)) and (layer0_outputs(7731)));
    layer1_outputs(2723) <= not(layer0_outputs(4731));
    layer1_outputs(2724) <= not(layer0_outputs(636));
    layer1_outputs(2725) <= not((layer0_outputs(2795)) or (layer0_outputs(25)));
    layer1_outputs(2726) <= layer0_outputs(5126);
    layer1_outputs(2727) <= layer0_outputs(5679);
    layer1_outputs(2728) <= not(layer0_outputs(6493)) or (layer0_outputs(8639));
    layer1_outputs(2729) <= (layer0_outputs(9068)) and not (layer0_outputs(9330));
    layer1_outputs(2730) <= layer0_outputs(9969);
    layer1_outputs(2731) <= not(layer0_outputs(6872)) or (layer0_outputs(7795));
    layer1_outputs(2732) <= not(layer0_outputs(2089));
    layer1_outputs(2733) <= (layer0_outputs(9991)) and not (layer0_outputs(8814));
    layer1_outputs(2734) <= not(layer0_outputs(6576));
    layer1_outputs(2735) <= not(layer0_outputs(6756));
    layer1_outputs(2736) <= not((layer0_outputs(4750)) and (layer0_outputs(3536)));
    layer1_outputs(2737) <= not(layer0_outputs(9031)) or (layer0_outputs(1830));
    layer1_outputs(2738) <= not(layer0_outputs(5406));
    layer1_outputs(2739) <= layer0_outputs(6483);
    layer1_outputs(2740) <= not((layer0_outputs(3344)) or (layer0_outputs(3181)));
    layer1_outputs(2741) <= layer0_outputs(6062);
    layer1_outputs(2742) <= layer0_outputs(7289);
    layer1_outputs(2743) <= not(layer0_outputs(6437));
    layer1_outputs(2744) <= '0';
    layer1_outputs(2745) <= (layer0_outputs(7383)) and not (layer0_outputs(4589));
    layer1_outputs(2746) <= not(layer0_outputs(7256));
    layer1_outputs(2747) <= not((layer0_outputs(3459)) xor (layer0_outputs(8315)));
    layer1_outputs(2748) <= (layer0_outputs(2427)) and not (layer0_outputs(7712));
    layer1_outputs(2749) <= layer0_outputs(4130);
    layer1_outputs(2750) <= not((layer0_outputs(6143)) or (layer0_outputs(3573)));
    layer1_outputs(2751) <= layer0_outputs(4318);
    layer1_outputs(2752) <= not(layer0_outputs(4644));
    layer1_outputs(2753) <= (layer0_outputs(4343)) and not (layer0_outputs(4106));
    layer1_outputs(2754) <= layer0_outputs(8289);
    layer1_outputs(2755) <= (layer0_outputs(6781)) or (layer0_outputs(10061));
    layer1_outputs(2756) <= not(layer0_outputs(8118));
    layer1_outputs(2757) <= (layer0_outputs(5626)) and not (layer0_outputs(337));
    layer1_outputs(2758) <= not(layer0_outputs(7025));
    layer1_outputs(2759) <= not(layer0_outputs(4359));
    layer1_outputs(2760) <= (layer0_outputs(1045)) and (layer0_outputs(778));
    layer1_outputs(2761) <= not(layer0_outputs(4442));
    layer1_outputs(2762) <= not((layer0_outputs(1826)) or (layer0_outputs(8484)));
    layer1_outputs(2763) <= not(layer0_outputs(4964));
    layer1_outputs(2764) <= layer0_outputs(6651);
    layer1_outputs(2765) <= not(layer0_outputs(7767));
    layer1_outputs(2766) <= not(layer0_outputs(6623));
    layer1_outputs(2767) <= layer0_outputs(3283);
    layer1_outputs(2768) <= not(layer0_outputs(5844));
    layer1_outputs(2769) <= not(layer0_outputs(4878)) or (layer0_outputs(9052));
    layer1_outputs(2770) <= not((layer0_outputs(5055)) or (layer0_outputs(3250)));
    layer1_outputs(2771) <= not(layer0_outputs(9447)) or (layer0_outputs(4614));
    layer1_outputs(2772) <= not((layer0_outputs(7473)) xor (layer0_outputs(2430)));
    layer1_outputs(2773) <= layer0_outputs(3140);
    layer1_outputs(2774) <= not((layer0_outputs(2718)) and (layer0_outputs(4474)));
    layer1_outputs(2775) <= (layer0_outputs(7588)) and not (layer0_outputs(9401));
    layer1_outputs(2776) <= (layer0_outputs(4010)) and not (layer0_outputs(460));
    layer1_outputs(2777) <= (layer0_outputs(7688)) and (layer0_outputs(809));
    layer1_outputs(2778) <= not((layer0_outputs(8637)) and (layer0_outputs(7645)));
    layer1_outputs(2779) <= not((layer0_outputs(2653)) xor (layer0_outputs(1778)));
    layer1_outputs(2780) <= not((layer0_outputs(8872)) xor (layer0_outputs(219)));
    layer1_outputs(2781) <= not((layer0_outputs(6178)) xor (layer0_outputs(4159)));
    layer1_outputs(2782) <= not(layer0_outputs(1121));
    layer1_outputs(2783) <= (layer0_outputs(2306)) or (layer0_outputs(7400));
    layer1_outputs(2784) <= not(layer0_outputs(4447)) or (layer0_outputs(3647));
    layer1_outputs(2785) <= not((layer0_outputs(2181)) xor (layer0_outputs(5969)));
    layer1_outputs(2786) <= '0';
    layer1_outputs(2787) <= layer0_outputs(5678);
    layer1_outputs(2788) <= not(layer0_outputs(7319));
    layer1_outputs(2789) <= (layer0_outputs(1166)) and not (layer0_outputs(9417));
    layer1_outputs(2790) <= (layer0_outputs(5550)) and not (layer0_outputs(3230));
    layer1_outputs(2791) <= not(layer0_outputs(4478));
    layer1_outputs(2792) <= not((layer0_outputs(8507)) and (layer0_outputs(1132)));
    layer1_outputs(2793) <= not(layer0_outputs(5549));
    layer1_outputs(2794) <= not((layer0_outputs(3947)) xor (layer0_outputs(3126)));
    layer1_outputs(2795) <= (layer0_outputs(3903)) xor (layer0_outputs(7910));
    layer1_outputs(2796) <= (layer0_outputs(9166)) xor (layer0_outputs(6641));
    layer1_outputs(2797) <= (layer0_outputs(6805)) xor (layer0_outputs(6714));
    layer1_outputs(2798) <= layer0_outputs(1383);
    layer1_outputs(2799) <= (layer0_outputs(7628)) xor (layer0_outputs(9611));
    layer1_outputs(2800) <= not(layer0_outputs(3667));
    layer1_outputs(2801) <= not((layer0_outputs(5346)) and (layer0_outputs(6444)));
    layer1_outputs(2802) <= not(layer0_outputs(1409));
    layer1_outputs(2803) <= not((layer0_outputs(3158)) xor (layer0_outputs(1192)));
    layer1_outputs(2804) <= not(layer0_outputs(5306)) or (layer0_outputs(6584));
    layer1_outputs(2805) <= (layer0_outputs(9875)) xor (layer0_outputs(4676));
    layer1_outputs(2806) <= layer0_outputs(5908);
    layer1_outputs(2807) <= (layer0_outputs(3214)) and not (layer0_outputs(8665));
    layer1_outputs(2808) <= (layer0_outputs(6678)) or (layer0_outputs(7509));
    layer1_outputs(2809) <= (layer0_outputs(1978)) and not (layer0_outputs(4756));
    layer1_outputs(2810) <= (layer0_outputs(992)) and not (layer0_outputs(7189));
    layer1_outputs(2811) <= (layer0_outputs(7618)) or (layer0_outputs(7323));
    layer1_outputs(2812) <= not(layer0_outputs(3267));
    layer1_outputs(2813) <= not(layer0_outputs(4868)) or (layer0_outputs(3469));
    layer1_outputs(2814) <= layer0_outputs(241);
    layer1_outputs(2815) <= layer0_outputs(6516);
    layer1_outputs(2816) <= not(layer0_outputs(8769)) or (layer0_outputs(5882));
    layer1_outputs(2817) <= (layer0_outputs(8287)) and not (layer0_outputs(8678));
    layer1_outputs(2818) <= (layer0_outputs(7332)) and not (layer0_outputs(8222));
    layer1_outputs(2819) <= '0';
    layer1_outputs(2820) <= (layer0_outputs(9888)) or (layer0_outputs(3447));
    layer1_outputs(2821) <= '1';
    layer1_outputs(2822) <= not((layer0_outputs(7003)) or (layer0_outputs(6334)));
    layer1_outputs(2823) <= layer0_outputs(93);
    layer1_outputs(2824) <= not((layer0_outputs(3753)) and (layer0_outputs(5267)));
    layer1_outputs(2825) <= not(layer0_outputs(1049)) or (layer0_outputs(314));
    layer1_outputs(2826) <= (layer0_outputs(6654)) and (layer0_outputs(4776));
    layer1_outputs(2827) <= (layer0_outputs(3692)) and (layer0_outputs(9500));
    layer1_outputs(2828) <= layer0_outputs(3589);
    layer1_outputs(2829) <= (layer0_outputs(7057)) or (layer0_outputs(9563));
    layer1_outputs(2830) <= layer0_outputs(219);
    layer1_outputs(2831) <= not(layer0_outputs(2147)) or (layer0_outputs(5876));
    layer1_outputs(2832) <= (layer0_outputs(3156)) and (layer0_outputs(6243));
    layer1_outputs(2833) <= layer0_outputs(2610);
    layer1_outputs(2834) <= not(layer0_outputs(4722)) or (layer0_outputs(8030));
    layer1_outputs(2835) <= (layer0_outputs(5217)) and not (layer0_outputs(6826));
    layer1_outputs(2836) <= not(layer0_outputs(2412)) or (layer0_outputs(4843));
    layer1_outputs(2837) <= not(layer0_outputs(175));
    layer1_outputs(2838) <= (layer0_outputs(5726)) xor (layer0_outputs(2760));
    layer1_outputs(2839) <= not(layer0_outputs(4015));
    layer1_outputs(2840) <= not((layer0_outputs(8726)) or (layer0_outputs(1086)));
    layer1_outputs(2841) <= layer0_outputs(1453);
    layer1_outputs(2842) <= not((layer0_outputs(7151)) and (layer0_outputs(6844)));
    layer1_outputs(2843) <= (layer0_outputs(113)) and not (layer0_outputs(7543));
    layer1_outputs(2844) <= not(layer0_outputs(1736));
    layer1_outputs(2845) <= layer0_outputs(4751);
    layer1_outputs(2846) <= (layer0_outputs(4951)) or (layer0_outputs(7831));
    layer1_outputs(2847) <= layer0_outputs(3721);
    layer1_outputs(2848) <= not(layer0_outputs(3824));
    layer1_outputs(2849) <= (layer0_outputs(5101)) xor (layer0_outputs(5197));
    layer1_outputs(2850) <= not(layer0_outputs(8328));
    layer1_outputs(2851) <= not((layer0_outputs(9636)) and (layer0_outputs(2870)));
    layer1_outputs(2852) <= (layer0_outputs(6241)) and (layer0_outputs(9399));
    layer1_outputs(2853) <= not(layer0_outputs(5078)) or (layer0_outputs(3306));
    layer1_outputs(2854) <= (layer0_outputs(10031)) and not (layer0_outputs(9123));
    layer1_outputs(2855) <= (layer0_outputs(6204)) and not (layer0_outputs(7707));
    layer1_outputs(2856) <= (layer0_outputs(1656)) and (layer0_outputs(2556));
    layer1_outputs(2857) <= layer0_outputs(8558);
    layer1_outputs(2858) <= (layer0_outputs(914)) xor (layer0_outputs(9609));
    layer1_outputs(2859) <= not((layer0_outputs(395)) and (layer0_outputs(3717)));
    layer1_outputs(2860) <= not(layer0_outputs(6968));
    layer1_outputs(2861) <= layer0_outputs(6467);
    layer1_outputs(2862) <= (layer0_outputs(4585)) and (layer0_outputs(619));
    layer1_outputs(2863) <= (layer0_outputs(398)) xor (layer0_outputs(5464));
    layer1_outputs(2864) <= not(layer0_outputs(1361)) or (layer0_outputs(2228));
    layer1_outputs(2865) <= (layer0_outputs(9853)) and not (layer0_outputs(9566));
    layer1_outputs(2866) <= (layer0_outputs(5954)) and not (layer0_outputs(8972));
    layer1_outputs(2867) <= (layer0_outputs(5601)) and not (layer0_outputs(6109));
    layer1_outputs(2868) <= not(layer0_outputs(9768)) or (layer0_outputs(2245));
    layer1_outputs(2869) <= layer0_outputs(4755);
    layer1_outputs(2870) <= not(layer0_outputs(3736)) or (layer0_outputs(7873));
    layer1_outputs(2871) <= (layer0_outputs(6130)) and (layer0_outputs(6640));
    layer1_outputs(2872) <= not(layer0_outputs(284));
    layer1_outputs(2873) <= layer0_outputs(5637);
    layer1_outputs(2874) <= not((layer0_outputs(2799)) and (layer0_outputs(6595)));
    layer1_outputs(2875) <= (layer0_outputs(8153)) and not (layer0_outputs(4425));
    layer1_outputs(2876) <= (layer0_outputs(6296)) xor (layer0_outputs(7168));
    layer1_outputs(2877) <= layer0_outputs(7642);
    layer1_outputs(2878) <= (layer0_outputs(6380)) and not (layer0_outputs(6197));
    layer1_outputs(2879) <= (layer0_outputs(1487)) and not (layer0_outputs(2958));
    layer1_outputs(2880) <= (layer0_outputs(958)) and not (layer0_outputs(3963));
    layer1_outputs(2881) <= layer0_outputs(2515);
    layer1_outputs(2882) <= (layer0_outputs(9161)) and (layer0_outputs(2893));
    layer1_outputs(2883) <= layer0_outputs(931);
    layer1_outputs(2884) <= not((layer0_outputs(4915)) or (layer0_outputs(3009)));
    layer1_outputs(2885) <= (layer0_outputs(9687)) or (layer0_outputs(6407));
    layer1_outputs(2886) <= layer0_outputs(614);
    layer1_outputs(2887) <= layer0_outputs(494);
    layer1_outputs(2888) <= not((layer0_outputs(7292)) and (layer0_outputs(8541)));
    layer1_outputs(2889) <= not((layer0_outputs(7013)) xor (layer0_outputs(8550)));
    layer1_outputs(2890) <= not(layer0_outputs(1714)) or (layer0_outputs(1534));
    layer1_outputs(2891) <= not(layer0_outputs(7754)) or (layer0_outputs(10149));
    layer1_outputs(2892) <= not(layer0_outputs(8803)) or (layer0_outputs(7257));
    layer1_outputs(2893) <= layer0_outputs(198);
    layer1_outputs(2894) <= (layer0_outputs(277)) and not (layer0_outputs(5215));
    layer1_outputs(2895) <= not((layer0_outputs(1074)) xor (layer0_outputs(1997)));
    layer1_outputs(2896) <= not(layer0_outputs(8924));
    layer1_outputs(2897) <= not((layer0_outputs(159)) xor (layer0_outputs(8438)));
    layer1_outputs(2898) <= not(layer0_outputs(885));
    layer1_outputs(2899) <= (layer0_outputs(2795)) and not (layer0_outputs(3717));
    layer1_outputs(2900) <= (layer0_outputs(8983)) and not (layer0_outputs(4543));
    layer1_outputs(2901) <= not((layer0_outputs(497)) and (layer0_outputs(2354)));
    layer1_outputs(2902) <= '1';
    layer1_outputs(2903) <= (layer0_outputs(1971)) and (layer0_outputs(5599));
    layer1_outputs(2904) <= not((layer0_outputs(5584)) or (layer0_outputs(1118)));
    layer1_outputs(2905) <= not((layer0_outputs(6985)) xor (layer0_outputs(3064)));
    layer1_outputs(2906) <= (layer0_outputs(1070)) and not (layer0_outputs(3921));
    layer1_outputs(2907) <= not(layer0_outputs(9129)) or (layer0_outputs(8690));
    layer1_outputs(2908) <= '0';
    layer1_outputs(2909) <= layer0_outputs(7674);
    layer1_outputs(2910) <= (layer0_outputs(362)) xor (layer0_outputs(4104));
    layer1_outputs(2911) <= not(layer0_outputs(9389)) or (layer0_outputs(3094));
    layer1_outputs(2912) <= not((layer0_outputs(491)) and (layer0_outputs(7091)));
    layer1_outputs(2913) <= (layer0_outputs(4775)) xor (layer0_outputs(5715));
    layer1_outputs(2914) <= (layer0_outputs(7697)) and (layer0_outputs(10203));
    layer1_outputs(2915) <= not(layer0_outputs(4012));
    layer1_outputs(2916) <= (layer0_outputs(2216)) and not (layer0_outputs(4967));
    layer1_outputs(2917) <= (layer0_outputs(4840)) xor (layer0_outputs(4339));
    layer1_outputs(2918) <= (layer0_outputs(124)) and not (layer0_outputs(6786));
    layer1_outputs(2919) <= not((layer0_outputs(7023)) xor (layer0_outputs(6012)));
    layer1_outputs(2920) <= not((layer0_outputs(4890)) xor (layer0_outputs(9673)));
    layer1_outputs(2921) <= not(layer0_outputs(9353));
    layer1_outputs(2922) <= not(layer0_outputs(9221)) or (layer0_outputs(9881));
    layer1_outputs(2923) <= layer0_outputs(7511);
    layer1_outputs(2924) <= not(layer0_outputs(3519));
    layer1_outputs(2925) <= not((layer0_outputs(6107)) and (layer0_outputs(3943)));
    layer1_outputs(2926) <= not((layer0_outputs(9543)) xor (layer0_outputs(7943)));
    layer1_outputs(2927) <= not((layer0_outputs(4900)) xor (layer0_outputs(238)));
    layer1_outputs(2928) <= (layer0_outputs(7639)) and not (layer0_outputs(5103));
    layer1_outputs(2929) <= not(layer0_outputs(9546)) or (layer0_outputs(6135));
    layer1_outputs(2930) <= layer0_outputs(2139);
    layer1_outputs(2931) <= not((layer0_outputs(7670)) or (layer0_outputs(7029)));
    layer1_outputs(2932) <= layer0_outputs(9047);
    layer1_outputs(2933) <= layer0_outputs(6355);
    layer1_outputs(2934) <= not(layer0_outputs(8342)) or (layer0_outputs(3803));
    layer1_outputs(2935) <= not(layer0_outputs(8860));
    layer1_outputs(2936) <= (layer0_outputs(5351)) xor (layer0_outputs(4372));
    layer1_outputs(2937) <= not(layer0_outputs(3134)) or (layer0_outputs(6815));
    layer1_outputs(2938) <= (layer0_outputs(2071)) and not (layer0_outputs(8391));
    layer1_outputs(2939) <= not(layer0_outputs(5628)) or (layer0_outputs(4391));
    layer1_outputs(2940) <= (layer0_outputs(4943)) and not (layer0_outputs(2763));
    layer1_outputs(2941) <= not(layer0_outputs(2387));
    layer1_outputs(2942) <= not(layer0_outputs(4116)) or (layer0_outputs(6688));
    layer1_outputs(2943) <= not(layer0_outputs(1894));
    layer1_outputs(2944) <= layer0_outputs(10093);
    layer1_outputs(2945) <= not(layer0_outputs(599));
    layer1_outputs(2946) <= (layer0_outputs(4700)) or (layer0_outputs(1371));
    layer1_outputs(2947) <= not((layer0_outputs(6809)) or (layer0_outputs(3979)));
    layer1_outputs(2948) <= layer0_outputs(9686);
    layer1_outputs(2949) <= (layer0_outputs(1948)) and not (layer0_outputs(7502));
    layer1_outputs(2950) <= (layer0_outputs(5670)) and not (layer0_outputs(840));
    layer1_outputs(2951) <= (layer0_outputs(3355)) and not (layer0_outputs(5439));
    layer1_outputs(2952) <= not(layer0_outputs(577));
    layer1_outputs(2953) <= not((layer0_outputs(6354)) xor (layer0_outputs(8407)));
    layer1_outputs(2954) <= not((layer0_outputs(716)) or (layer0_outputs(8190)));
    layer1_outputs(2955) <= layer0_outputs(7378);
    layer1_outputs(2956) <= not(layer0_outputs(3168));
    layer1_outputs(2957) <= layer0_outputs(2213);
    layer1_outputs(2958) <= not(layer0_outputs(6698));
    layer1_outputs(2959) <= (layer0_outputs(8266)) and not (layer0_outputs(4357));
    layer1_outputs(2960) <= (layer0_outputs(631)) or (layer0_outputs(2771));
    layer1_outputs(2961) <= not((layer0_outputs(5075)) or (layer0_outputs(5814)));
    layer1_outputs(2962) <= layer0_outputs(8681);
    layer1_outputs(2963) <= (layer0_outputs(7800)) and not (layer0_outputs(2917));
    layer1_outputs(2964) <= not(layer0_outputs(1399));
    layer1_outputs(2965) <= (layer0_outputs(8302)) and not (layer0_outputs(1584));
    layer1_outputs(2966) <= not(layer0_outputs(8124));
    layer1_outputs(2967) <= layer0_outputs(3549);
    layer1_outputs(2968) <= (layer0_outputs(8333)) or (layer0_outputs(4967));
    layer1_outputs(2969) <= layer0_outputs(4842);
    layer1_outputs(2970) <= not((layer0_outputs(3480)) xor (layer0_outputs(6170)));
    layer1_outputs(2971) <= not((layer0_outputs(1057)) or (layer0_outputs(6544)));
    layer1_outputs(2972) <= (layer0_outputs(833)) xor (layer0_outputs(1955));
    layer1_outputs(2973) <= not((layer0_outputs(3956)) or (layer0_outputs(4438)));
    layer1_outputs(2974) <= (layer0_outputs(8240)) xor (layer0_outputs(7563));
    layer1_outputs(2975) <= layer0_outputs(5369);
    layer1_outputs(2976) <= not((layer0_outputs(5462)) xor (layer0_outputs(6778)));
    layer1_outputs(2977) <= (layer0_outputs(8943)) and not (layer0_outputs(1615));
    layer1_outputs(2978) <= not(layer0_outputs(3608));
    layer1_outputs(2979) <= not(layer0_outputs(9587));
    layer1_outputs(2980) <= not((layer0_outputs(1224)) xor (layer0_outputs(4870)));
    layer1_outputs(2981) <= not(layer0_outputs(5128)) or (layer0_outputs(3855));
    layer1_outputs(2982) <= not(layer0_outputs(2858)) or (layer0_outputs(672));
    layer1_outputs(2983) <= layer0_outputs(10126);
    layer1_outputs(2984) <= not(layer0_outputs(8060));
    layer1_outputs(2985) <= not(layer0_outputs(5733));
    layer1_outputs(2986) <= not(layer0_outputs(6804)) or (layer0_outputs(2975));
    layer1_outputs(2987) <= not((layer0_outputs(4867)) and (layer0_outputs(10190)));
    layer1_outputs(2988) <= (layer0_outputs(5718)) or (layer0_outputs(8993));
    layer1_outputs(2989) <= layer0_outputs(2468);
    layer1_outputs(2990) <= not(layer0_outputs(4059));
    layer1_outputs(2991) <= not((layer0_outputs(9785)) and (layer0_outputs(4404)));
    layer1_outputs(2992) <= not((layer0_outputs(1831)) or (layer0_outputs(115)));
    layer1_outputs(2993) <= not((layer0_outputs(8250)) and (layer0_outputs(3171)));
    layer1_outputs(2994) <= (layer0_outputs(1884)) and not (layer0_outputs(6849));
    layer1_outputs(2995) <= not(layer0_outputs(9545));
    layer1_outputs(2996) <= (layer0_outputs(130)) and (layer0_outputs(4474));
    layer1_outputs(2997) <= not((layer0_outputs(3130)) or (layer0_outputs(6850)));
    layer1_outputs(2998) <= layer0_outputs(6736);
    layer1_outputs(2999) <= not(layer0_outputs(7492)) or (layer0_outputs(2347));
    layer1_outputs(3000) <= (layer0_outputs(995)) and (layer0_outputs(8368));
    layer1_outputs(3001) <= (layer0_outputs(3852)) and not (layer0_outputs(8100));
    layer1_outputs(3002) <= not(layer0_outputs(3229));
    layer1_outputs(3003) <= layer0_outputs(2701);
    layer1_outputs(3004) <= (layer0_outputs(8084)) or (layer0_outputs(10084));
    layer1_outputs(3005) <= not((layer0_outputs(5214)) or (layer0_outputs(6784)));
    layer1_outputs(3006) <= not(layer0_outputs(4618));
    layer1_outputs(3007) <= not(layer0_outputs(215)) or (layer0_outputs(10231));
    layer1_outputs(3008) <= not(layer0_outputs(424)) or (layer0_outputs(7443));
    layer1_outputs(3009) <= not(layer0_outputs(1175)) or (layer0_outputs(1695));
    layer1_outputs(3010) <= layer0_outputs(8603);
    layer1_outputs(3011) <= not(layer0_outputs(7405));
    layer1_outputs(3012) <= not(layer0_outputs(381));
    layer1_outputs(3013) <= not((layer0_outputs(8820)) xor (layer0_outputs(215)));
    layer1_outputs(3014) <= not((layer0_outputs(8168)) xor (layer0_outputs(799)));
    layer1_outputs(3015) <= not((layer0_outputs(5034)) and (layer0_outputs(9552)));
    layer1_outputs(3016) <= (layer0_outputs(490)) and (layer0_outputs(7927));
    layer1_outputs(3017) <= (layer0_outputs(5784)) xor (layer0_outputs(4096));
    layer1_outputs(3018) <= not(layer0_outputs(4720));
    layer1_outputs(3019) <= (layer0_outputs(7390)) and not (layer0_outputs(3749));
    layer1_outputs(3020) <= not(layer0_outputs(4324));
    layer1_outputs(3021) <= (layer0_outputs(10190)) xor (layer0_outputs(3326));
    layer1_outputs(3022) <= not(layer0_outputs(4634)) or (layer0_outputs(1232));
    layer1_outputs(3023) <= not(layer0_outputs(333)) or (layer0_outputs(4642));
    layer1_outputs(3024) <= (layer0_outputs(9279)) and not (layer0_outputs(7376));
    layer1_outputs(3025) <= (layer0_outputs(45)) xor (layer0_outputs(10106));
    layer1_outputs(3026) <= (layer0_outputs(10043)) and not (layer0_outputs(2847));
    layer1_outputs(3027) <= (layer0_outputs(3585)) and (layer0_outputs(582));
    layer1_outputs(3028) <= not(layer0_outputs(8106)) or (layer0_outputs(6827));
    layer1_outputs(3029) <= not(layer0_outputs(5538)) or (layer0_outputs(2359));
    layer1_outputs(3030) <= (layer0_outputs(1014)) xor (layer0_outputs(3152));
    layer1_outputs(3031) <= (layer0_outputs(4754)) and not (layer0_outputs(9988));
    layer1_outputs(3032) <= (layer0_outputs(1591)) and not (layer0_outputs(6603));
    layer1_outputs(3033) <= (layer0_outputs(44)) and not (layer0_outputs(3450));
    layer1_outputs(3034) <= '1';
    layer1_outputs(3035) <= (layer0_outputs(5912)) xor (layer0_outputs(363));
    layer1_outputs(3036) <= (layer0_outputs(4792)) xor (layer0_outputs(9271));
    layer1_outputs(3037) <= not(layer0_outputs(5557));
    layer1_outputs(3038) <= not(layer0_outputs(4669)) or (layer0_outputs(7436));
    layer1_outputs(3039) <= (layer0_outputs(2122)) and (layer0_outputs(2995));
    layer1_outputs(3040) <= not((layer0_outputs(9690)) and (layer0_outputs(443)));
    layer1_outputs(3041) <= (layer0_outputs(3604)) xor (layer0_outputs(2044));
    layer1_outputs(3042) <= not(layer0_outputs(8101));
    layer1_outputs(3043) <= layer0_outputs(803);
    layer1_outputs(3044) <= not(layer0_outputs(2895)) or (layer0_outputs(6541));
    layer1_outputs(3045) <= not(layer0_outputs(2948));
    layer1_outputs(3046) <= layer0_outputs(6408);
    layer1_outputs(3047) <= (layer0_outputs(9129)) and not (layer0_outputs(9458));
    layer1_outputs(3048) <= not((layer0_outputs(5247)) and (layer0_outputs(7043)));
    layer1_outputs(3049) <= (layer0_outputs(3989)) or (layer0_outputs(8128));
    layer1_outputs(3050) <= layer0_outputs(1685);
    layer1_outputs(3051) <= not(layer0_outputs(8863));
    layer1_outputs(3052) <= not((layer0_outputs(5052)) or (layer0_outputs(2675)));
    layer1_outputs(3053) <= not((layer0_outputs(3971)) and (layer0_outputs(4945)));
    layer1_outputs(3054) <= (layer0_outputs(1621)) xor (layer0_outputs(5072));
    layer1_outputs(3055) <= not(layer0_outputs(3010));
    layer1_outputs(3056) <= not((layer0_outputs(9190)) and (layer0_outputs(5426)));
    layer1_outputs(3057) <= (layer0_outputs(8243)) or (layer0_outputs(1840));
    layer1_outputs(3058) <= '0';
    layer1_outputs(3059) <= not(layer0_outputs(6828));
    layer1_outputs(3060) <= (layer0_outputs(1526)) and not (layer0_outputs(4578));
    layer1_outputs(3061) <= '1';
    layer1_outputs(3062) <= not(layer0_outputs(2574)) or (layer0_outputs(9014));
    layer1_outputs(3063) <= not((layer0_outputs(8747)) and (layer0_outputs(113)));
    layer1_outputs(3064) <= not((layer0_outputs(9966)) or (layer0_outputs(2113)));
    layer1_outputs(3065) <= '0';
    layer1_outputs(3066) <= (layer0_outputs(9562)) and not (layer0_outputs(2819));
    layer1_outputs(3067) <= (layer0_outputs(6441)) and not (layer0_outputs(1868));
    layer1_outputs(3068) <= (layer0_outputs(5136)) and (layer0_outputs(9244));
    layer1_outputs(3069) <= not((layer0_outputs(9409)) and (layer0_outputs(1502)));
    layer1_outputs(3070) <= not(layer0_outputs(6377)) or (layer0_outputs(7637));
    layer1_outputs(3071) <= layer0_outputs(5066);
    layer1_outputs(3072) <= not((layer0_outputs(682)) xor (layer0_outputs(4590)));
    layer1_outputs(3073) <= (layer0_outputs(1630)) and not (layer0_outputs(8257));
    layer1_outputs(3074) <= (layer0_outputs(6002)) and not (layer0_outputs(248));
    layer1_outputs(3075) <= not((layer0_outputs(8775)) and (layer0_outputs(8970)));
    layer1_outputs(3076) <= not((layer0_outputs(9857)) or (layer0_outputs(3067)));
    layer1_outputs(3077) <= not(layer0_outputs(8258));
    layer1_outputs(3078) <= (layer0_outputs(4477)) or (layer0_outputs(7741));
    layer1_outputs(3079) <= not(layer0_outputs(9753)) or (layer0_outputs(9505));
    layer1_outputs(3080) <= layer0_outputs(5666);
    layer1_outputs(3081) <= layer0_outputs(9850);
    layer1_outputs(3082) <= layer0_outputs(782);
    layer1_outputs(3083) <= layer0_outputs(7019);
    layer1_outputs(3084) <= not(layer0_outputs(4018));
    layer1_outputs(3085) <= not(layer0_outputs(4088)) or (layer0_outputs(4264));
    layer1_outputs(3086) <= layer0_outputs(3368);
    layer1_outputs(3087) <= (layer0_outputs(4491)) and (layer0_outputs(1699));
    layer1_outputs(3088) <= not(layer0_outputs(6619)) or (layer0_outputs(5118));
    layer1_outputs(3089) <= not((layer0_outputs(3384)) or (layer0_outputs(9806)));
    layer1_outputs(3090) <= not(layer0_outputs(2699)) or (layer0_outputs(2340));
    layer1_outputs(3091) <= not(layer0_outputs(4427)) or (layer0_outputs(2429));
    layer1_outputs(3092) <= (layer0_outputs(7584)) and (layer0_outputs(5026));
    layer1_outputs(3093) <= not(layer0_outputs(3603));
    layer1_outputs(3094) <= not(layer0_outputs(5338));
    layer1_outputs(3095) <= layer0_outputs(4836);
    layer1_outputs(3096) <= (layer0_outputs(1243)) xor (layer0_outputs(1717));
    layer1_outputs(3097) <= '1';
    layer1_outputs(3098) <= layer0_outputs(6819);
    layer1_outputs(3099) <= not(layer0_outputs(2882)) or (layer0_outputs(6319));
    layer1_outputs(3100) <= not(layer0_outputs(9450));
    layer1_outputs(3101) <= not(layer0_outputs(2856));
    layer1_outputs(3102) <= not(layer0_outputs(4161)) or (layer0_outputs(746));
    layer1_outputs(3103) <= layer0_outputs(8731);
    layer1_outputs(3104) <= layer0_outputs(2943);
    layer1_outputs(3105) <= (layer0_outputs(4152)) and (layer0_outputs(6996));
    layer1_outputs(3106) <= not(layer0_outputs(2384)) or (layer0_outputs(8318));
    layer1_outputs(3107) <= not(layer0_outputs(9283)) or (layer0_outputs(6172));
    layer1_outputs(3108) <= not(layer0_outputs(6206)) or (layer0_outputs(3320));
    layer1_outputs(3109) <= layer0_outputs(8406);
    layer1_outputs(3110) <= (layer0_outputs(3262)) and (layer0_outputs(5508));
    layer1_outputs(3111) <= (layer0_outputs(9708)) and not (layer0_outputs(9314));
    layer1_outputs(3112) <= layer0_outputs(9926);
    layer1_outputs(3113) <= not((layer0_outputs(1934)) and (layer0_outputs(9579)));
    layer1_outputs(3114) <= layer0_outputs(4753);
    layer1_outputs(3115) <= layer0_outputs(9337);
    layer1_outputs(3116) <= (layer0_outputs(5150)) and not (layer0_outputs(2418));
    layer1_outputs(3117) <= not(layer0_outputs(4535)) or (layer0_outputs(5667));
    layer1_outputs(3118) <= layer0_outputs(7284);
    layer1_outputs(3119) <= '0';
    layer1_outputs(3120) <= not(layer0_outputs(3075));
    layer1_outputs(3121) <= (layer0_outputs(10111)) and not (layer0_outputs(1538));
    layer1_outputs(3122) <= layer0_outputs(9712);
    layer1_outputs(3123) <= not(layer0_outputs(4593));
    layer1_outputs(3124) <= (layer0_outputs(5645)) and not (layer0_outputs(7851));
    layer1_outputs(3125) <= not(layer0_outputs(3114)) or (layer0_outputs(2746));
    layer1_outputs(3126) <= not((layer0_outputs(6481)) or (layer0_outputs(6574)));
    layer1_outputs(3127) <= not(layer0_outputs(7333));
    layer1_outputs(3128) <= not(layer0_outputs(3244));
    layer1_outputs(3129) <= layer0_outputs(6475);
    layer1_outputs(3130) <= layer0_outputs(2902);
    layer1_outputs(3131) <= not((layer0_outputs(3937)) and (layer0_outputs(5345)));
    layer1_outputs(3132) <= not(layer0_outputs(6694));
    layer1_outputs(3133) <= not(layer0_outputs(5559));
    layer1_outputs(3134) <= not(layer0_outputs(4181));
    layer1_outputs(3135) <= (layer0_outputs(4264)) and not (layer0_outputs(5080));
    layer1_outputs(3136) <= not(layer0_outputs(3846)) or (layer0_outputs(5495));
    layer1_outputs(3137) <= layer0_outputs(4583);
    layer1_outputs(3138) <= not((layer0_outputs(1227)) and (layer0_outputs(4932)));
    layer1_outputs(3139) <= (layer0_outputs(7194)) or (layer0_outputs(2128));
    layer1_outputs(3140) <= (layer0_outputs(652)) and not (layer0_outputs(192));
    layer1_outputs(3141) <= not(layer0_outputs(3131));
    layer1_outputs(3142) <= not(layer0_outputs(7232)) or (layer0_outputs(5504));
    layer1_outputs(3143) <= layer0_outputs(4431);
    layer1_outputs(3144) <= layer0_outputs(10056);
    layer1_outputs(3145) <= (layer0_outputs(3433)) and (layer0_outputs(5165));
    layer1_outputs(3146) <= layer0_outputs(4559);
    layer1_outputs(3147) <= layer0_outputs(4573);
    layer1_outputs(3148) <= not(layer0_outputs(1776)) or (layer0_outputs(4176));
    layer1_outputs(3149) <= not(layer0_outputs(5697)) or (layer0_outputs(8741));
    layer1_outputs(3150) <= not((layer0_outputs(7583)) or (layer0_outputs(1739)));
    layer1_outputs(3151) <= (layer0_outputs(6379)) and not (layer0_outputs(3028));
    layer1_outputs(3152) <= (layer0_outputs(2869)) and (layer0_outputs(9205));
    layer1_outputs(3153) <= (layer0_outputs(8859)) and (layer0_outputs(275));
    layer1_outputs(3154) <= (layer0_outputs(9188)) and (layer0_outputs(8729));
    layer1_outputs(3155) <= layer0_outputs(3336);
    layer1_outputs(3156) <= (layer0_outputs(2816)) or (layer0_outputs(1593));
    layer1_outputs(3157) <= not(layer0_outputs(1610));
    layer1_outputs(3158) <= not((layer0_outputs(5148)) and (layer0_outputs(6711)));
    layer1_outputs(3159) <= layer0_outputs(3246);
    layer1_outputs(3160) <= not(layer0_outputs(1064)) or (layer0_outputs(2677));
    layer1_outputs(3161) <= not(layer0_outputs(10047));
    layer1_outputs(3162) <= layer0_outputs(823);
    layer1_outputs(3163) <= (layer0_outputs(6645)) or (layer0_outputs(5244));
    layer1_outputs(3164) <= not(layer0_outputs(5220));
    layer1_outputs(3165) <= not(layer0_outputs(1696));
    layer1_outputs(3166) <= (layer0_outputs(5749)) xor (layer0_outputs(7279));
    layer1_outputs(3167) <= not(layer0_outputs(8524));
    layer1_outputs(3168) <= not(layer0_outputs(4281)) or (layer0_outputs(9237));
    layer1_outputs(3169) <= not((layer0_outputs(3223)) or (layer0_outputs(8851)));
    layer1_outputs(3170) <= not((layer0_outputs(3671)) xor (layer0_outputs(3531)));
    layer1_outputs(3171) <= not(layer0_outputs(5255));
    layer1_outputs(3172) <= not(layer0_outputs(4719));
    layer1_outputs(3173) <= not((layer0_outputs(7014)) or (layer0_outputs(10087)));
    layer1_outputs(3174) <= not(layer0_outputs(6787));
    layer1_outputs(3175) <= not(layer0_outputs(2542));
    layer1_outputs(3176) <= layer0_outputs(4100);
    layer1_outputs(3177) <= (layer0_outputs(632)) and not (layer0_outputs(8197));
    layer1_outputs(3178) <= not(layer0_outputs(5447));
    layer1_outputs(3179) <= (layer0_outputs(333)) and (layer0_outputs(6059));
    layer1_outputs(3180) <= (layer0_outputs(5980)) or (layer0_outputs(3170));
    layer1_outputs(3181) <= (layer0_outputs(10120)) xor (layer0_outputs(4556));
    layer1_outputs(3182) <= (layer0_outputs(10160)) and (layer0_outputs(7673));
    layer1_outputs(3183) <= (layer0_outputs(6916)) and not (layer0_outputs(5337));
    layer1_outputs(3184) <= layer0_outputs(8013);
    layer1_outputs(3185) <= not(layer0_outputs(4914));
    layer1_outputs(3186) <= layer0_outputs(8165);
    layer1_outputs(3187) <= (layer0_outputs(9006)) and not (layer0_outputs(6564));
    layer1_outputs(3188) <= '0';
    layer1_outputs(3189) <= layer0_outputs(9962);
    layer1_outputs(3190) <= (layer0_outputs(9253)) and not (layer0_outputs(2792));
    layer1_outputs(3191) <= not((layer0_outputs(674)) and (layer0_outputs(8916)));
    layer1_outputs(3192) <= (layer0_outputs(5490)) and (layer0_outputs(6056));
    layer1_outputs(3193) <= not(layer0_outputs(1120));
    layer1_outputs(3194) <= layer0_outputs(3048);
    layer1_outputs(3195) <= layer0_outputs(4805);
    layer1_outputs(3196) <= (layer0_outputs(1414)) and (layer0_outputs(6994));
    layer1_outputs(3197) <= layer0_outputs(6171);
    layer1_outputs(3198) <= layer0_outputs(10029);
    layer1_outputs(3199) <= not((layer0_outputs(7334)) and (layer0_outputs(8569)));
    layer1_outputs(3200) <= not(layer0_outputs(5151)) or (layer0_outputs(9940));
    layer1_outputs(3201) <= layer0_outputs(3431);
    layer1_outputs(3202) <= not((layer0_outputs(440)) and (layer0_outputs(9944)));
    layer1_outputs(3203) <= '0';
    layer1_outputs(3204) <= not(layer0_outputs(1000));
    layer1_outputs(3205) <= not(layer0_outputs(3149)) or (layer0_outputs(2088));
    layer1_outputs(3206) <= (layer0_outputs(2539)) xor (layer0_outputs(603));
    layer1_outputs(3207) <= not((layer0_outputs(5942)) or (layer0_outputs(6690)));
    layer1_outputs(3208) <= (layer0_outputs(9347)) or (layer0_outputs(5479));
    layer1_outputs(3209) <= not(layer0_outputs(9913)) or (layer0_outputs(9942));
    layer1_outputs(3210) <= (layer0_outputs(3987)) and not (layer0_outputs(5424));
    layer1_outputs(3211) <= (layer0_outputs(123)) and not (layer0_outputs(3256));
    layer1_outputs(3212) <= layer0_outputs(3108);
    layer1_outputs(3213) <= (layer0_outputs(7542)) and not (layer0_outputs(8113));
    layer1_outputs(3214) <= not((layer0_outputs(1423)) or (layer0_outputs(2054)));
    layer1_outputs(3215) <= not(layer0_outputs(9730)) or (layer0_outputs(8005));
    layer1_outputs(3216) <= layer0_outputs(4047);
    layer1_outputs(3217) <= not(layer0_outputs(8839)) or (layer0_outputs(1076));
    layer1_outputs(3218) <= (layer0_outputs(8752)) xor (layer0_outputs(2531));
    layer1_outputs(3219) <= not(layer0_outputs(610));
    layer1_outputs(3220) <= not((layer0_outputs(7596)) or (layer0_outputs(1140)));
    layer1_outputs(3221) <= not((layer0_outputs(2652)) or (layer0_outputs(9692)));
    layer1_outputs(3222) <= '0';
    layer1_outputs(3223) <= layer0_outputs(10208);
    layer1_outputs(3224) <= not((layer0_outputs(10125)) xor (layer0_outputs(6289)));
    layer1_outputs(3225) <= not((layer0_outputs(7280)) or (layer0_outputs(3239)));
    layer1_outputs(3226) <= layer0_outputs(4603);
    layer1_outputs(3227) <= layer0_outputs(6669);
    layer1_outputs(3228) <= not(layer0_outputs(8828)) or (layer0_outputs(734));
    layer1_outputs(3229) <= not(layer0_outputs(5283)) or (layer0_outputs(3568));
    layer1_outputs(3230) <= (layer0_outputs(965)) and not (layer0_outputs(8316));
    layer1_outputs(3231) <= not(layer0_outputs(8994));
    layer1_outputs(3232) <= not(layer0_outputs(7093)) or (layer0_outputs(3558));
    layer1_outputs(3233) <= not(layer0_outputs(3867));
    layer1_outputs(3234) <= (layer0_outputs(621)) and not (layer0_outputs(4210));
    layer1_outputs(3235) <= not(layer0_outputs(4178));
    layer1_outputs(3236) <= (layer0_outputs(6982)) or (layer0_outputs(9101));
    layer1_outputs(3237) <= not(layer0_outputs(3133));
    layer1_outputs(3238) <= not((layer0_outputs(8361)) or (layer0_outputs(3808)));
    layer1_outputs(3239) <= not(layer0_outputs(3057));
    layer1_outputs(3240) <= layer0_outputs(7562);
    layer1_outputs(3241) <= not(layer0_outputs(3845));
    layer1_outputs(3242) <= not(layer0_outputs(7085)) or (layer0_outputs(4169));
    layer1_outputs(3243) <= (layer0_outputs(363)) and not (layer0_outputs(1247));
    layer1_outputs(3244) <= (layer0_outputs(8000)) and not (layer0_outputs(2939));
    layer1_outputs(3245) <= not(layer0_outputs(5603)) or (layer0_outputs(209));
    layer1_outputs(3246) <= (layer0_outputs(4686)) and not (layer0_outputs(1020));
    layer1_outputs(3247) <= not(layer0_outputs(5287)) or (layer0_outputs(9985));
    layer1_outputs(3248) <= not(layer0_outputs(607));
    layer1_outputs(3249) <= not(layer0_outputs(5252)) or (layer0_outputs(3476));
    layer1_outputs(3250) <= not(layer0_outputs(1729));
    layer1_outputs(3251) <= (layer0_outputs(2714)) and not (layer0_outputs(3881));
    layer1_outputs(3252) <= (layer0_outputs(1095)) xor (layer0_outputs(9067));
    layer1_outputs(3253) <= not((layer0_outputs(5501)) or (layer0_outputs(4921)));
    layer1_outputs(3254) <= layer0_outputs(6567);
    layer1_outputs(3255) <= not((layer0_outputs(2021)) and (layer0_outputs(2228)));
    layer1_outputs(3256) <= (layer0_outputs(6712)) or (layer0_outputs(874));
    layer1_outputs(3257) <= (layer0_outputs(5678)) and not (layer0_outputs(5236));
    layer1_outputs(3258) <= not(layer0_outputs(3134)) or (layer0_outputs(8083));
    layer1_outputs(3259) <= not(layer0_outputs(9613)) or (layer0_outputs(2190));
    layer1_outputs(3260) <= not((layer0_outputs(5513)) or (layer0_outputs(5310)));
    layer1_outputs(3261) <= not((layer0_outputs(3865)) and (layer0_outputs(9788)));
    layer1_outputs(3262) <= layer0_outputs(4917);
    layer1_outputs(3263) <= not((layer0_outputs(3748)) and (layer0_outputs(5494)));
    layer1_outputs(3264) <= not(layer0_outputs(6378)) or (layer0_outputs(5265));
    layer1_outputs(3265) <= not((layer0_outputs(660)) and (layer0_outputs(4840)));
    layer1_outputs(3266) <= (layer0_outputs(3466)) and not (layer0_outputs(6886));
    layer1_outputs(3267) <= (layer0_outputs(6573)) xor (layer0_outputs(9582));
    layer1_outputs(3268) <= (layer0_outputs(8186)) and not (layer0_outputs(8312));
    layer1_outputs(3269) <= not(layer0_outputs(7380));
    layer1_outputs(3270) <= layer0_outputs(8826);
    layer1_outputs(3271) <= layer0_outputs(8248);
    layer1_outputs(3272) <= not(layer0_outputs(5700));
    layer1_outputs(3273) <= (layer0_outputs(343)) xor (layer0_outputs(1129));
    layer1_outputs(3274) <= not(layer0_outputs(3678));
    layer1_outputs(3275) <= not(layer0_outputs(6834));
    layer1_outputs(3276) <= (layer0_outputs(1250)) and (layer0_outputs(8570));
    layer1_outputs(3277) <= not(layer0_outputs(126)) or (layer0_outputs(5234));
    layer1_outputs(3278) <= not(layer0_outputs(7438));
    layer1_outputs(3279) <= layer0_outputs(5090);
    layer1_outputs(3280) <= (layer0_outputs(718)) or (layer0_outputs(3766));
    layer1_outputs(3281) <= not((layer0_outputs(10227)) xor (layer0_outputs(762)));
    layer1_outputs(3282) <= layer0_outputs(9152);
    layer1_outputs(3283) <= (layer0_outputs(1643)) xor (layer0_outputs(3157));
    layer1_outputs(3284) <= not(layer0_outputs(3967));
    layer1_outputs(3285) <= layer0_outputs(6205);
    layer1_outputs(3286) <= not(layer0_outputs(8964));
    layer1_outputs(3287) <= (layer0_outputs(870)) or (layer0_outputs(4670));
    layer1_outputs(3288) <= '0';
    layer1_outputs(3289) <= (layer0_outputs(8948)) and not (layer0_outputs(3164));
    layer1_outputs(3290) <= not((layer0_outputs(6035)) and (layer0_outputs(1961)));
    layer1_outputs(3291) <= not((layer0_outputs(4676)) xor (layer0_outputs(3617)));
    layer1_outputs(3292) <= not(layer0_outputs(10171)) or (layer0_outputs(3622));
    layer1_outputs(3293) <= not((layer0_outputs(7071)) or (layer0_outputs(1639)));
    layer1_outputs(3294) <= layer0_outputs(1459);
    layer1_outputs(3295) <= layer0_outputs(2445);
    layer1_outputs(3296) <= layer0_outputs(8646);
    layer1_outputs(3297) <= not(layer0_outputs(357)) or (layer0_outputs(2385));
    layer1_outputs(3298) <= (layer0_outputs(8309)) xor (layer0_outputs(9035));
    layer1_outputs(3299) <= (layer0_outputs(668)) and not (layer0_outputs(1464));
    layer1_outputs(3300) <= layer0_outputs(150);
    layer1_outputs(3301) <= not(layer0_outputs(9357)) or (layer0_outputs(2151));
    layer1_outputs(3302) <= not((layer0_outputs(7595)) xor (layer0_outputs(4325)));
    layer1_outputs(3303) <= not((layer0_outputs(1829)) or (layer0_outputs(1924)));
    layer1_outputs(3304) <= layer0_outputs(3793);
    layer1_outputs(3305) <= not((layer0_outputs(3992)) xor (layer0_outputs(4374)));
    layer1_outputs(3306) <= not(layer0_outputs(7847));
    layer1_outputs(3307) <= not(layer0_outputs(7069));
    layer1_outputs(3308) <= (layer0_outputs(9003)) or (layer0_outputs(8091));
    layer1_outputs(3309) <= layer0_outputs(10006);
    layer1_outputs(3310) <= (layer0_outputs(1049)) and not (layer0_outputs(9887));
    layer1_outputs(3311) <= not(layer0_outputs(490));
    layer1_outputs(3312) <= not(layer0_outputs(4606));
    layer1_outputs(3313) <= (layer0_outputs(3434)) and not (layer0_outputs(1386));
    layer1_outputs(3314) <= not(layer0_outputs(7187));
    layer1_outputs(3315) <= layer0_outputs(9283);
    layer1_outputs(3316) <= not((layer0_outputs(781)) or (layer0_outputs(3605)));
    layer1_outputs(3317) <= layer0_outputs(3088);
    layer1_outputs(3318) <= (layer0_outputs(2334)) and not (layer0_outputs(1910));
    layer1_outputs(3319) <= (layer0_outputs(819)) xor (layer0_outputs(6458));
    layer1_outputs(3320) <= not((layer0_outputs(2422)) xor (layer0_outputs(3645)));
    layer1_outputs(3321) <= not(layer0_outputs(7480));
    layer1_outputs(3322) <= not(layer0_outputs(9571)) or (layer0_outputs(5581));
    layer1_outputs(3323) <= not(layer0_outputs(9681)) or (layer0_outputs(8320));
    layer1_outputs(3324) <= not(layer0_outputs(2929)) or (layer0_outputs(8147));
    layer1_outputs(3325) <= not((layer0_outputs(2437)) or (layer0_outputs(5566)));
    layer1_outputs(3326) <= not((layer0_outputs(6633)) xor (layer0_outputs(4107)));
    layer1_outputs(3327) <= layer0_outputs(1644);
    layer1_outputs(3328) <= layer0_outputs(272);
    layer1_outputs(3329) <= not(layer0_outputs(3919)) or (layer0_outputs(8579));
    layer1_outputs(3330) <= not((layer0_outputs(2373)) xor (layer0_outputs(9779)));
    layer1_outputs(3331) <= not(layer0_outputs(5857)) or (layer0_outputs(1678));
    layer1_outputs(3332) <= (layer0_outputs(6)) or (layer0_outputs(4089));
    layer1_outputs(3333) <= not(layer0_outputs(1717));
    layer1_outputs(3334) <= layer0_outputs(9465);
    layer1_outputs(3335) <= not((layer0_outputs(5233)) and (layer0_outputs(3783)));
    layer1_outputs(3336) <= not(layer0_outputs(10221)) or (layer0_outputs(7246));
    layer1_outputs(3337) <= not(layer0_outputs(2981)) or (layer0_outputs(4697));
    layer1_outputs(3338) <= not(layer0_outputs(6591));
    layer1_outputs(3339) <= (layer0_outputs(7109)) and not (layer0_outputs(8278));
    layer1_outputs(3340) <= (layer0_outputs(8778)) and not (layer0_outputs(4201));
    layer1_outputs(3341) <= '0';
    layer1_outputs(3342) <= not(layer0_outputs(2014));
    layer1_outputs(3343) <= not(layer0_outputs(5482)) or (layer0_outputs(931));
    layer1_outputs(3344) <= (layer0_outputs(7967)) and (layer0_outputs(2018));
    layer1_outputs(3345) <= (layer0_outputs(679)) and not (layer0_outputs(10026));
    layer1_outputs(3346) <= layer0_outputs(2339);
    layer1_outputs(3347) <= layer0_outputs(3470);
    layer1_outputs(3348) <= (layer0_outputs(4550)) and (layer0_outputs(2621));
    layer1_outputs(3349) <= (layer0_outputs(1018)) and (layer0_outputs(2432));
    layer1_outputs(3350) <= not(layer0_outputs(9724)) or (layer0_outputs(573));
    layer1_outputs(3351) <= (layer0_outputs(4217)) and (layer0_outputs(86));
    layer1_outputs(3352) <= not(layer0_outputs(8897));
    layer1_outputs(3353) <= not(layer0_outputs(8456));
    layer1_outputs(3354) <= (layer0_outputs(6436)) xor (layer0_outputs(100));
    layer1_outputs(3355) <= not(layer0_outputs(8779));
    layer1_outputs(3356) <= not(layer0_outputs(300));
    layer1_outputs(3357) <= (layer0_outputs(5446)) and not (layer0_outputs(5521));
    layer1_outputs(3358) <= not(layer0_outputs(8399));
    layer1_outputs(3359) <= '0';
    layer1_outputs(3360) <= not(layer0_outputs(5356));
    layer1_outputs(3361) <= (layer0_outputs(1391)) and not (layer0_outputs(7150));
    layer1_outputs(3362) <= layer0_outputs(8883);
    layer1_outputs(3363) <= not((layer0_outputs(5385)) or (layer0_outputs(5870)));
    layer1_outputs(3364) <= not(layer0_outputs(2163));
    layer1_outputs(3365) <= (layer0_outputs(2470)) and not (layer0_outputs(7059));
    layer1_outputs(3366) <= (layer0_outputs(5790)) and not (layer0_outputs(9391));
    layer1_outputs(3367) <= not(layer0_outputs(9195));
    layer1_outputs(3368) <= not(layer0_outputs(2618));
    layer1_outputs(3369) <= layer0_outputs(5071);
    layer1_outputs(3370) <= layer0_outputs(9841);
    layer1_outputs(3371) <= not((layer0_outputs(9559)) xor (layer0_outputs(1154)));
    layer1_outputs(3372) <= not((layer0_outputs(2985)) and (layer0_outputs(9893)));
    layer1_outputs(3373) <= not(layer0_outputs(8074)) or (layer0_outputs(10158));
    layer1_outputs(3374) <= '0';
    layer1_outputs(3375) <= layer0_outputs(506);
    layer1_outputs(3376) <= not(layer0_outputs(7983));
    layer1_outputs(3377) <= not(layer0_outputs(1763)) or (layer0_outputs(7487));
    layer1_outputs(3378) <= (layer0_outputs(2841)) or (layer0_outputs(6387));
    layer1_outputs(3379) <= '1';
    layer1_outputs(3380) <= (layer0_outputs(8986)) xor (layer0_outputs(4628));
    layer1_outputs(3381) <= (layer0_outputs(262)) and not (layer0_outputs(995));
    layer1_outputs(3382) <= not((layer0_outputs(4842)) and (layer0_outputs(6705)));
    layer1_outputs(3383) <= layer0_outputs(10151);
    layer1_outputs(3384) <= not(layer0_outputs(4280));
    layer1_outputs(3385) <= not(layer0_outputs(971));
    layer1_outputs(3386) <= layer0_outputs(10009);
    layer1_outputs(3387) <= layer0_outputs(8039);
    layer1_outputs(3388) <= (layer0_outputs(3098)) or (layer0_outputs(10083));
    layer1_outputs(3389) <= (layer0_outputs(3020)) and not (layer0_outputs(2572));
    layer1_outputs(3390) <= layer0_outputs(8901);
    layer1_outputs(3391) <= not((layer0_outputs(8348)) and (layer0_outputs(2509)));
    layer1_outputs(3392) <= (layer0_outputs(9949)) and (layer0_outputs(8160));
    layer1_outputs(3393) <= not((layer0_outputs(9817)) or (layer0_outputs(2109)));
    layer1_outputs(3394) <= layer0_outputs(2765);
    layer1_outputs(3395) <= layer0_outputs(9044);
    layer1_outputs(3396) <= layer0_outputs(5365);
    layer1_outputs(3397) <= not(layer0_outputs(2433));
    layer1_outputs(3398) <= not(layer0_outputs(3719));
    layer1_outputs(3399) <= layer0_outputs(533);
    layer1_outputs(3400) <= not((layer0_outputs(10183)) or (layer0_outputs(3851)));
    layer1_outputs(3401) <= not((layer0_outputs(1030)) or (layer0_outputs(9177)));
    layer1_outputs(3402) <= not(layer0_outputs(10164));
    layer1_outputs(3403) <= not(layer0_outputs(5918));
    layer1_outputs(3404) <= not(layer0_outputs(5675));
    layer1_outputs(3405) <= layer0_outputs(4780);
    layer1_outputs(3406) <= '1';
    layer1_outputs(3407) <= layer0_outputs(10068);
    layer1_outputs(3408) <= layer0_outputs(3525);
    layer1_outputs(3409) <= (layer0_outputs(1667)) and not (layer0_outputs(6339));
    layer1_outputs(3410) <= not(layer0_outputs(669)) or (layer0_outputs(3897));
    layer1_outputs(3411) <= not((layer0_outputs(7965)) and (layer0_outputs(5375)));
    layer1_outputs(3412) <= (layer0_outputs(917)) and not (layer0_outputs(2952));
    layer1_outputs(3413) <= not(layer0_outputs(7860)) or (layer0_outputs(5092));
    layer1_outputs(3414) <= layer0_outputs(1291);
    layer1_outputs(3415) <= layer0_outputs(6733);
    layer1_outputs(3416) <= not(layer0_outputs(9007));
    layer1_outputs(3417) <= not((layer0_outputs(8992)) or (layer0_outputs(1571)));
    layer1_outputs(3418) <= not(layer0_outputs(998));
    layer1_outputs(3419) <= not(layer0_outputs(2507));
    layer1_outputs(3420) <= (layer0_outputs(4368)) or (layer0_outputs(8309));
    layer1_outputs(3421) <= (layer0_outputs(8600)) and (layer0_outputs(2218));
    layer1_outputs(3422) <= (layer0_outputs(8985)) and (layer0_outputs(8239));
    layer1_outputs(3423) <= layer0_outputs(6893);
    layer1_outputs(3424) <= (layer0_outputs(7377)) and not (layer0_outputs(3176));
    layer1_outputs(3425) <= not((layer0_outputs(5060)) xor (layer0_outputs(5627)));
    layer1_outputs(3426) <= not((layer0_outputs(3432)) or (layer0_outputs(9772)));
    layer1_outputs(3427) <= (layer0_outputs(5420)) or (layer0_outputs(644));
    layer1_outputs(3428) <= (layer0_outputs(300)) and (layer0_outputs(4675));
    layer1_outputs(3429) <= not((layer0_outputs(1184)) or (layer0_outputs(5441)));
    layer1_outputs(3430) <= not((layer0_outputs(292)) and (layer0_outputs(5525)));
    layer1_outputs(3431) <= not((layer0_outputs(9781)) xor (layer0_outputs(10140)));
    layer1_outputs(3432) <= layer0_outputs(10033);
    layer1_outputs(3433) <= (layer0_outputs(5325)) and not (layer0_outputs(3986));
    layer1_outputs(3434) <= '1';
    layer1_outputs(3435) <= not(layer0_outputs(2366)) or (layer0_outputs(7733));
    layer1_outputs(3436) <= layer0_outputs(7554);
    layer1_outputs(3437) <= (layer0_outputs(7932)) and not (layer0_outputs(2185));
    layer1_outputs(3438) <= layer0_outputs(9367);
    layer1_outputs(3439) <= (layer0_outputs(7444)) xor (layer0_outputs(8688));
    layer1_outputs(3440) <= not(layer0_outputs(7721)) or (layer0_outputs(2595));
    layer1_outputs(3441) <= not(layer0_outputs(3893));
    layer1_outputs(3442) <= not(layer0_outputs(9705));
    layer1_outputs(3443) <= not(layer0_outputs(5941));
    layer1_outputs(3444) <= not(layer0_outputs(1732));
    layer1_outputs(3445) <= (layer0_outputs(5251)) xor (layer0_outputs(5434));
    layer1_outputs(3446) <= not(layer0_outputs(7521)) or (layer0_outputs(7585));
    layer1_outputs(3447) <= not(layer0_outputs(1399));
    layer1_outputs(3448) <= (layer0_outputs(5688)) xor (layer0_outputs(4197));
    layer1_outputs(3449) <= (layer0_outputs(8198)) and not (layer0_outputs(10045));
    layer1_outputs(3450) <= not((layer0_outputs(6513)) xor (layer0_outputs(2528)));
    layer1_outputs(3451) <= (layer0_outputs(4846)) xor (layer0_outputs(6475));
    layer1_outputs(3452) <= layer0_outputs(2079);
    layer1_outputs(3453) <= not((layer0_outputs(5113)) xor (layer0_outputs(9019)));
    layer1_outputs(3454) <= not((layer0_outputs(1748)) and (layer0_outputs(2772)));
    layer1_outputs(3455) <= not(layer0_outputs(2503)) or (layer0_outputs(1914));
    layer1_outputs(3456) <= not(layer0_outputs(2035));
    layer1_outputs(3457) <= (layer0_outputs(2345)) and not (layer0_outputs(8352));
    layer1_outputs(3458) <= layer0_outputs(2226);
    layer1_outputs(3459) <= not(layer0_outputs(10215)) or (layer0_outputs(3621));
    layer1_outputs(3460) <= not(layer0_outputs(9675)) or (layer0_outputs(5428));
    layer1_outputs(3461) <= not(layer0_outputs(6573));
    layer1_outputs(3462) <= (layer0_outputs(8354)) and (layer0_outputs(4982));
    layer1_outputs(3463) <= (layer0_outputs(1150)) and (layer0_outputs(8704));
    layer1_outputs(3464) <= (layer0_outputs(5759)) and not (layer0_outputs(479));
    layer1_outputs(3465) <= (layer0_outputs(3705)) and not (layer0_outputs(1898));
    layer1_outputs(3466) <= not(layer0_outputs(3810)) or (layer0_outputs(1663));
    layer1_outputs(3467) <= not(layer0_outputs(3970));
    layer1_outputs(3468) <= (layer0_outputs(6292)) and (layer0_outputs(5147));
    layer1_outputs(3469) <= (layer0_outputs(7937)) or (layer0_outputs(7035));
    layer1_outputs(3470) <= (layer0_outputs(178)) or (layer0_outputs(9586));
    layer1_outputs(3471) <= (layer0_outputs(5702)) and not (layer0_outputs(2921));
    layer1_outputs(3472) <= not(layer0_outputs(9010));
    layer1_outputs(3473) <= (layer0_outputs(9553)) and (layer0_outputs(1141));
    layer1_outputs(3474) <= (layer0_outputs(7059)) or (layer0_outputs(1587));
    layer1_outputs(3475) <= not(layer0_outputs(8642));
    layer1_outputs(3476) <= not((layer0_outputs(6718)) xor (layer0_outputs(7144)));
    layer1_outputs(3477) <= not(layer0_outputs(1936));
    layer1_outputs(3478) <= (layer0_outputs(690)) and not (layer0_outputs(1384));
    layer1_outputs(3479) <= '1';
    layer1_outputs(3480) <= not(layer0_outputs(5961));
    layer1_outputs(3481) <= layer0_outputs(3152);
    layer1_outputs(3482) <= not((layer0_outputs(991)) or (layer0_outputs(277)));
    layer1_outputs(3483) <= (layer0_outputs(568)) and (layer0_outputs(3995));
    layer1_outputs(3484) <= not((layer0_outputs(367)) or (layer0_outputs(6741)));
    layer1_outputs(3485) <= not((layer0_outputs(3546)) or (layer0_outputs(9953)));
    layer1_outputs(3486) <= (layer0_outputs(8732)) and not (layer0_outputs(4081));
    layer1_outputs(3487) <= (layer0_outputs(8412)) and (layer0_outputs(7598));
    layer1_outputs(3488) <= not(layer0_outputs(10134));
    layer1_outputs(3489) <= layer0_outputs(8662);
    layer1_outputs(3490) <= not(layer0_outputs(2766)) or (layer0_outputs(9426));
    layer1_outputs(3491) <= not(layer0_outputs(10107)) or (layer0_outputs(2442));
    layer1_outputs(3492) <= layer0_outputs(4101);
    layer1_outputs(3493) <= not(layer0_outputs(5786)) or (layer0_outputs(4392));
    layer1_outputs(3494) <= '1';
    layer1_outputs(3495) <= (layer0_outputs(9346)) and not (layer0_outputs(2382));
    layer1_outputs(3496) <= not(layer0_outputs(3368));
    layer1_outputs(3497) <= not(layer0_outputs(3006)) or (layer0_outputs(6015));
    layer1_outputs(3498) <= not((layer0_outputs(3194)) and (layer0_outputs(6875)));
    layer1_outputs(3499) <= layer0_outputs(4612);
    layer1_outputs(3500) <= not(layer0_outputs(404));
    layer1_outputs(3501) <= (layer0_outputs(1395)) or (layer0_outputs(874));
    layer1_outputs(3502) <= not((layer0_outputs(2720)) xor (layer0_outputs(7734)));
    layer1_outputs(3503) <= not((layer0_outputs(883)) or (layer0_outputs(9985)));
    layer1_outputs(3504) <= not((layer0_outputs(3132)) or (layer0_outputs(4216)));
    layer1_outputs(3505) <= layer0_outputs(7992);
    layer1_outputs(3506) <= not(layer0_outputs(4108)) or (layer0_outputs(4553));
    layer1_outputs(3507) <= layer0_outputs(7812);
    layer1_outputs(3508) <= (layer0_outputs(2294)) and (layer0_outputs(17));
    layer1_outputs(3509) <= (layer0_outputs(1524)) and (layer0_outputs(3554));
    layer1_outputs(3510) <= (layer0_outputs(2842)) and not (layer0_outputs(8942));
    layer1_outputs(3511) <= not(layer0_outputs(2179)) or (layer0_outputs(847));
    layer1_outputs(3512) <= (layer0_outputs(904)) or (layer0_outputs(301));
    layer1_outputs(3513) <= not(layer0_outputs(8373));
    layer1_outputs(3514) <= not(layer0_outputs(10114)) or (layer0_outputs(2604));
    layer1_outputs(3515) <= not((layer0_outputs(8025)) or (layer0_outputs(8580)));
    layer1_outputs(3516) <= layer0_outputs(3446);
    layer1_outputs(3517) <= not(layer0_outputs(125));
    layer1_outputs(3518) <= (layer0_outputs(8687)) and not (layer0_outputs(2206));
    layer1_outputs(3519) <= layer0_outputs(9581);
    layer1_outputs(3520) <= not(layer0_outputs(1949));
    layer1_outputs(3521) <= (layer0_outputs(1465)) xor (layer0_outputs(9285));
    layer1_outputs(3522) <= not(layer0_outputs(10106));
    layer1_outputs(3523) <= layer0_outputs(7702);
    layer1_outputs(3524) <= not(layer0_outputs(8221));
    layer1_outputs(3525) <= not((layer0_outputs(9430)) xor (layer0_outputs(3453)));
    layer1_outputs(3526) <= not((layer0_outputs(4021)) xor (layer0_outputs(9948)));
    layer1_outputs(3527) <= layer0_outputs(2741);
    layer1_outputs(3528) <= (layer0_outputs(2899)) or (layer0_outputs(9834));
    layer1_outputs(3529) <= (layer0_outputs(8144)) xor (layer0_outputs(9687));
    layer1_outputs(3530) <= (layer0_outputs(6354)) or (layer0_outputs(5146));
    layer1_outputs(3531) <= (layer0_outputs(5218)) and not (layer0_outputs(445));
    layer1_outputs(3532) <= not(layer0_outputs(1203));
    layer1_outputs(3533) <= (layer0_outputs(1823)) and not (layer0_outputs(3454));
    layer1_outputs(3534) <= not(layer0_outputs(3278));
    layer1_outputs(3535) <= not(layer0_outputs(5510));
    layer1_outputs(3536) <= (layer0_outputs(1145)) or (layer0_outputs(7835));
    layer1_outputs(3537) <= (layer0_outputs(9519)) or (layer0_outputs(8536));
    layer1_outputs(3538) <= not(layer0_outputs(9585)) or (layer0_outputs(8544));
    layer1_outputs(3539) <= (layer0_outputs(5413)) and not (layer0_outputs(5445));
    layer1_outputs(3540) <= not(layer0_outputs(3098));
    layer1_outputs(3541) <= not(layer0_outputs(9108));
    layer1_outputs(3542) <= '0';
    layer1_outputs(3543) <= not(layer0_outputs(8534)) or (layer0_outputs(9245));
    layer1_outputs(3544) <= not(layer0_outputs(9470));
    layer1_outputs(3545) <= (layer0_outputs(8385)) and (layer0_outputs(6746));
    layer1_outputs(3546) <= not(layer0_outputs(4370));
    layer1_outputs(3547) <= (layer0_outputs(5622)) and not (layer0_outputs(3951));
    layer1_outputs(3548) <= (layer0_outputs(2949)) xor (layer0_outputs(8275));
    layer1_outputs(3549) <= not(layer0_outputs(8556));
    layer1_outputs(3550) <= not(layer0_outputs(3085)) or (layer0_outputs(7147));
    layer1_outputs(3551) <= not(layer0_outputs(8636));
    layer1_outputs(3552) <= (layer0_outputs(9529)) and not (layer0_outputs(2926));
    layer1_outputs(3553) <= not(layer0_outputs(6756));
    layer1_outputs(3554) <= layer0_outputs(4350);
    layer1_outputs(3555) <= not(layer0_outputs(3917));
    layer1_outputs(3556) <= (layer0_outputs(274)) and (layer0_outputs(6930));
    layer1_outputs(3557) <= not(layer0_outputs(8009));
    layer1_outputs(3558) <= not(layer0_outputs(7593));
    layer1_outputs(3559) <= layer0_outputs(5657);
    layer1_outputs(3560) <= layer0_outputs(356);
    layer1_outputs(3561) <= layer0_outputs(496);
    layer1_outputs(3562) <= (layer0_outputs(8037)) or (layer0_outputs(9491));
    layer1_outputs(3563) <= layer0_outputs(3179);
    layer1_outputs(3564) <= not(layer0_outputs(1664));
    layer1_outputs(3565) <= not((layer0_outputs(4228)) and (layer0_outputs(9068)));
    layer1_outputs(3566) <= (layer0_outputs(4065)) and not (layer0_outputs(3437));
    layer1_outputs(3567) <= not(layer0_outputs(6037)) or (layer0_outputs(1807));
    layer1_outputs(3568) <= layer0_outputs(10233);
    layer1_outputs(3569) <= not((layer0_outputs(8735)) or (layer0_outputs(2344)));
    layer1_outputs(3570) <= (layer0_outputs(625)) and not (layer0_outputs(9845));
    layer1_outputs(3571) <= layer0_outputs(5730);
    layer1_outputs(3572) <= (layer0_outputs(3397)) xor (layer0_outputs(3441));
    layer1_outputs(3573) <= layer0_outputs(3568);
    layer1_outputs(3574) <= not((layer0_outputs(10198)) and (layer0_outputs(337)));
    layer1_outputs(3575) <= layer0_outputs(6471);
    layer1_outputs(3576) <= not(layer0_outputs(610));
    layer1_outputs(3577) <= not((layer0_outputs(4880)) or (layer0_outputs(195)));
    layer1_outputs(3578) <= layer0_outputs(6028);
    layer1_outputs(3579) <= (layer0_outputs(9083)) and not (layer0_outputs(9807));
    layer1_outputs(3580) <= not(layer0_outputs(9752)) or (layer0_outputs(981));
    layer1_outputs(3581) <= not(layer0_outputs(2157));
    layer1_outputs(3582) <= (layer0_outputs(1512)) or (layer0_outputs(7727));
    layer1_outputs(3583) <= layer0_outputs(6717);
    layer1_outputs(3584) <= not((layer0_outputs(471)) xor (layer0_outputs(6853)));
    layer1_outputs(3585) <= not(layer0_outputs(7083));
    layer1_outputs(3586) <= not(layer0_outputs(1756)) or (layer0_outputs(5481));
    layer1_outputs(3587) <= (layer0_outputs(2253)) and not (layer0_outputs(5700));
    layer1_outputs(3588) <= (layer0_outputs(132)) xor (layer0_outputs(4707));
    layer1_outputs(3589) <= layer0_outputs(6764);
    layer1_outputs(3590) <= not(layer0_outputs(1770)) or (layer0_outputs(3768));
    layer1_outputs(3591) <= not(layer0_outputs(9660));
    layer1_outputs(3592) <= not(layer0_outputs(6922)) or (layer0_outputs(3611));
    layer1_outputs(3593) <= layer0_outputs(7218);
    layer1_outputs(3594) <= '0';
    layer1_outputs(3595) <= layer0_outputs(677);
    layer1_outputs(3596) <= not((layer0_outputs(6689)) and (layer0_outputs(754)));
    layer1_outputs(3597) <= not((layer0_outputs(8548)) or (layer0_outputs(6133)));
    layer1_outputs(3598) <= layer0_outputs(3513);
    layer1_outputs(3599) <= layer0_outputs(9827);
    layer1_outputs(3600) <= not((layer0_outputs(1179)) and (layer0_outputs(2970)));
    layer1_outputs(3601) <= (layer0_outputs(2396)) xor (layer0_outputs(6157));
    layer1_outputs(3602) <= not((layer0_outputs(8459)) and (layer0_outputs(7049)));
    layer1_outputs(3603) <= not(layer0_outputs(4659)) or (layer0_outputs(1471));
    layer1_outputs(3604) <= not((layer0_outputs(6780)) or (layer0_outputs(4491)));
    layer1_outputs(3605) <= (layer0_outputs(3633)) and not (layer0_outputs(4481));
    layer1_outputs(3606) <= (layer0_outputs(2407)) and not (layer0_outputs(1845));
    layer1_outputs(3607) <= not(layer0_outputs(2670));
    layer1_outputs(3608) <= (layer0_outputs(725)) or (layer0_outputs(1364));
    layer1_outputs(3609) <= not(layer0_outputs(9199));
    layer1_outputs(3610) <= (layer0_outputs(4276)) or (layer0_outputs(10146));
    layer1_outputs(3611) <= not((layer0_outputs(7882)) xor (layer0_outputs(7194)));
    layer1_outputs(3612) <= (layer0_outputs(7770)) or (layer0_outputs(8799));
    layer1_outputs(3613) <= layer0_outputs(7713);
    layer1_outputs(3614) <= not(layer0_outputs(2101)) or (layer0_outputs(6269));
    layer1_outputs(3615) <= not(layer0_outputs(876)) or (layer0_outputs(5390));
    layer1_outputs(3616) <= not(layer0_outputs(4770));
    layer1_outputs(3617) <= (layer0_outputs(9794)) and (layer0_outputs(5673));
    layer1_outputs(3618) <= not(layer0_outputs(9890));
    layer1_outputs(3619) <= not((layer0_outputs(7307)) and (layer0_outputs(5326)));
    layer1_outputs(3620) <= (layer0_outputs(4075)) xor (layer0_outputs(1412));
    layer1_outputs(3621) <= (layer0_outputs(203)) and not (layer0_outputs(6770));
    layer1_outputs(3622) <= not((layer0_outputs(2814)) and (layer0_outputs(9778)));
    layer1_outputs(3623) <= not(layer0_outputs(5677)) or (layer0_outputs(458));
    layer1_outputs(3624) <= (layer0_outputs(7979)) or (layer0_outputs(8987));
    layer1_outputs(3625) <= not(layer0_outputs(600));
    layer1_outputs(3626) <= not(layer0_outputs(5057));
    layer1_outputs(3627) <= layer0_outputs(10003);
    layer1_outputs(3628) <= layer0_outputs(7407);
    layer1_outputs(3629) <= (layer0_outputs(2673)) and not (layer0_outputs(6260));
    layer1_outputs(3630) <= not((layer0_outputs(3685)) xor (layer0_outputs(1301)));
    layer1_outputs(3631) <= (layer0_outputs(7086)) and not (layer0_outputs(5076));
    layer1_outputs(3632) <= not(layer0_outputs(8314));
    layer1_outputs(3633) <= not(layer0_outputs(4432));
    layer1_outputs(3634) <= not(layer0_outputs(4228)) or (layer0_outputs(977));
    layer1_outputs(3635) <= (layer0_outputs(8227)) and not (layer0_outputs(5553));
    layer1_outputs(3636) <= layer0_outputs(5093);
    layer1_outputs(3637) <= not((layer0_outputs(8825)) and (layer0_outputs(1444)));
    layer1_outputs(3638) <= not((layer0_outputs(470)) and (layer0_outputs(2203)));
    layer1_outputs(3639) <= (layer0_outputs(1079)) and (layer0_outputs(879));
    layer1_outputs(3640) <= (layer0_outputs(1426)) or (layer0_outputs(3183));
    layer1_outputs(3641) <= (layer0_outputs(2807)) and not (layer0_outputs(8555));
    layer1_outputs(3642) <= (layer0_outputs(3306)) or (layer0_outputs(10093));
    layer1_outputs(3643) <= (layer0_outputs(5909)) or (layer0_outputs(3146));
    layer1_outputs(3644) <= (layer0_outputs(1738)) xor (layer0_outputs(2417));
    layer1_outputs(3645) <= not(layer0_outputs(781)) or (layer0_outputs(2731));
    layer1_outputs(3646) <= layer0_outputs(8287);
    layer1_outputs(3647) <= layer0_outputs(4698);
    layer1_outputs(3648) <= not((layer0_outputs(6169)) xor (layer0_outputs(5558)));
    layer1_outputs(3649) <= layer0_outputs(9622);
    layer1_outputs(3650) <= not(layer0_outputs(3064));
    layer1_outputs(3651) <= not(layer0_outputs(1374));
    layer1_outputs(3652) <= (layer0_outputs(10191)) or (layer0_outputs(3291));
    layer1_outputs(3653) <= layer0_outputs(482);
    layer1_outputs(3654) <= not(layer0_outputs(1316));
    layer1_outputs(3655) <= not(layer0_outputs(8268));
    layer1_outputs(3656) <= layer0_outputs(8720);
    layer1_outputs(3657) <= not((layer0_outputs(6337)) and (layer0_outputs(4850)));
    layer1_outputs(3658) <= not(layer0_outputs(9795)) or (layer0_outputs(9293));
    layer1_outputs(3659) <= layer0_outputs(6966);
    layer1_outputs(3660) <= not((layer0_outputs(3841)) or (layer0_outputs(9897)));
    layer1_outputs(3661) <= (layer0_outputs(8143)) and not (layer0_outputs(419));
    layer1_outputs(3662) <= (layer0_outputs(9258)) or (layer0_outputs(6284));
    layer1_outputs(3663) <= not(layer0_outputs(4265));
    layer1_outputs(3664) <= not(layer0_outputs(1873));
    layer1_outputs(3665) <= layer0_outputs(3304);
    layer1_outputs(3666) <= '1';
    layer1_outputs(3667) <= not(layer0_outputs(3865)) or (layer0_outputs(5605));
    layer1_outputs(3668) <= layer0_outputs(1726);
    layer1_outputs(3669) <= (layer0_outputs(8204)) or (layer0_outputs(1959));
    layer1_outputs(3670) <= not(layer0_outputs(4401)) or (layer0_outputs(3377));
    layer1_outputs(3671) <= layer0_outputs(2941);
    layer1_outputs(3672) <= layer0_outputs(10206);
    layer1_outputs(3673) <= not(layer0_outputs(1141));
    layer1_outputs(3674) <= not((layer0_outputs(1359)) xor (layer0_outputs(2415)));
    layer1_outputs(3675) <= not((layer0_outputs(8127)) xor (layer0_outputs(6798)));
    layer1_outputs(3676) <= not(layer0_outputs(6667));
    layer1_outputs(3677) <= not(layer0_outputs(10025));
    layer1_outputs(3678) <= (layer0_outputs(4783)) and not (layer0_outputs(9493));
    layer1_outputs(3679) <= not(layer0_outputs(4143));
    layer1_outputs(3680) <= layer0_outputs(2096);
    layer1_outputs(3681) <= (layer0_outputs(4029)) and not (layer0_outputs(9843));
    layer1_outputs(3682) <= (layer0_outputs(666)) xor (layer0_outputs(2862));
    layer1_outputs(3683) <= not((layer0_outputs(4171)) and (layer0_outputs(9397)));
    layer1_outputs(3684) <= (layer0_outputs(1782)) or (layer0_outputs(1945));
    layer1_outputs(3685) <= (layer0_outputs(1096)) and not (layer0_outputs(8958));
    layer1_outputs(3686) <= not((layer0_outputs(5027)) or (layer0_outputs(2267)));
    layer1_outputs(3687) <= not((layer0_outputs(5668)) or (layer0_outputs(6540)));
    layer1_outputs(3688) <= layer0_outputs(2754);
    layer1_outputs(3689) <= not((layer0_outputs(8893)) and (layer0_outputs(4118)));
    layer1_outputs(3690) <= (layer0_outputs(967)) and not (layer0_outputs(4886));
    layer1_outputs(3691) <= not(layer0_outputs(7300)) or (layer0_outputs(2045));
    layer1_outputs(3692) <= not((layer0_outputs(365)) xor (layer0_outputs(5980)));
    layer1_outputs(3693) <= not((layer0_outputs(9289)) and (layer0_outputs(6640)));
    layer1_outputs(3694) <= not(layer0_outputs(8413)) or (layer0_outputs(8467));
    layer1_outputs(3695) <= not(layer0_outputs(2060));
    layer1_outputs(3696) <= not((layer0_outputs(6689)) and (layer0_outputs(6310)));
    layer1_outputs(3697) <= not(layer0_outputs(1755)) or (layer0_outputs(9578));
    layer1_outputs(3698) <= (layer0_outputs(2629)) and not (layer0_outputs(7094));
    layer1_outputs(3699) <= (layer0_outputs(6552)) and not (layer0_outputs(6829));
    layer1_outputs(3700) <= not((layer0_outputs(9671)) or (layer0_outputs(901)));
    layer1_outputs(3701) <= not(layer0_outputs(6774)) or (layer0_outputs(7890));
    layer1_outputs(3702) <= layer0_outputs(9807);
    layer1_outputs(3703) <= (layer0_outputs(8096)) xor (layer0_outputs(2717));
    layer1_outputs(3704) <= (layer0_outputs(8132)) and not (layer0_outputs(2440));
    layer1_outputs(3705) <= layer0_outputs(9425);
    layer1_outputs(3706) <= (layer0_outputs(4171)) xor (layer0_outputs(3944));
    layer1_outputs(3707) <= (layer0_outputs(8118)) and not (layer0_outputs(3089));
    layer1_outputs(3708) <= (layer0_outputs(10100)) xor (layer0_outputs(3275));
    layer1_outputs(3709) <= layer0_outputs(4033);
    layer1_outputs(3710) <= '0';
    layer1_outputs(3711) <= (layer0_outputs(1787)) and not (layer0_outputs(10174));
    layer1_outputs(3712) <= not((layer0_outputs(9586)) xor (layer0_outputs(7515)));
    layer1_outputs(3713) <= (layer0_outputs(466)) and not (layer0_outputs(1285));
    layer1_outputs(3714) <= not(layer0_outputs(2669));
    layer1_outputs(3715) <= not(layer0_outputs(8081));
    layer1_outputs(3716) <= not(layer0_outputs(7122)) or (layer0_outputs(5911));
    layer1_outputs(3717) <= (layer0_outputs(9057)) or (layer0_outputs(1965));
    layer1_outputs(3718) <= not((layer0_outputs(3365)) or (layer0_outputs(6176)));
    layer1_outputs(3719) <= not((layer0_outputs(9989)) and (layer0_outputs(1)));
    layer1_outputs(3720) <= not(layer0_outputs(2103)) or (layer0_outputs(6048));
    layer1_outputs(3721) <= (layer0_outputs(6512)) xor (layer0_outputs(9671));
    layer1_outputs(3722) <= (layer0_outputs(4075)) and not (layer0_outputs(2963));
    layer1_outputs(3723) <= (layer0_outputs(8092)) or (layer0_outputs(2102));
    layer1_outputs(3724) <= '1';
    layer1_outputs(3725) <= not(layer0_outputs(10102));
    layer1_outputs(3726) <= not(layer0_outputs(4396)) or (layer0_outputs(338));
    layer1_outputs(3727) <= layer0_outputs(796);
    layer1_outputs(3728) <= not(layer0_outputs(6877));
    layer1_outputs(3729) <= layer0_outputs(1730);
    layer1_outputs(3730) <= not(layer0_outputs(5717));
    layer1_outputs(3731) <= not(layer0_outputs(2924)) or (layer0_outputs(10176));
    layer1_outputs(3732) <= not(layer0_outputs(221));
    layer1_outputs(3733) <= not(layer0_outputs(8397)) or (layer0_outputs(2575));
    layer1_outputs(3734) <= layer0_outputs(413);
    layer1_outputs(3735) <= (layer0_outputs(6115)) and not (layer0_outputs(69));
    layer1_outputs(3736) <= not(layer0_outputs(1568));
    layer1_outputs(3737) <= layer0_outputs(3634);
    layer1_outputs(3738) <= not(layer0_outputs(6620)) or (layer0_outputs(1852));
    layer1_outputs(3739) <= layer0_outputs(2015);
    layer1_outputs(3740) <= not((layer0_outputs(2055)) or (layer0_outputs(6115)));
    layer1_outputs(3741) <= not(layer0_outputs(1509));
    layer1_outputs(3742) <= layer0_outputs(4563);
    layer1_outputs(3743) <= (layer0_outputs(2036)) and not (layer0_outputs(10161));
    layer1_outputs(3744) <= not((layer0_outputs(2961)) xor (layer0_outputs(4193)));
    layer1_outputs(3745) <= (layer0_outputs(3370)) or (layer0_outputs(5249));
    layer1_outputs(3746) <= (layer0_outputs(422)) or (layer0_outputs(7274));
    layer1_outputs(3747) <= not(layer0_outputs(524));
    layer1_outputs(3748) <= layer0_outputs(5164);
    layer1_outputs(3749) <= (layer0_outputs(9299)) and not (layer0_outputs(2773));
    layer1_outputs(3750) <= not((layer0_outputs(6399)) or (layer0_outputs(4844)));
    layer1_outputs(3751) <= not(layer0_outputs(8729));
    layer1_outputs(3752) <= layer0_outputs(929);
    layer1_outputs(3753) <= layer0_outputs(6157);
    layer1_outputs(3754) <= layer0_outputs(4983);
    layer1_outputs(3755) <= not((layer0_outputs(8577)) or (layer0_outputs(8961)));
    layer1_outputs(3756) <= (layer0_outputs(8751)) or (layer0_outputs(8259));
    layer1_outputs(3757) <= not((layer0_outputs(7889)) or (layer0_outputs(3452)));
    layer1_outputs(3758) <= (layer0_outputs(6988)) and (layer0_outputs(2230));
    layer1_outputs(3759) <= not(layer0_outputs(8955));
    layer1_outputs(3760) <= not(layer0_outputs(5029));
    layer1_outputs(3761) <= not(layer0_outputs(4160));
    layer1_outputs(3762) <= layer0_outputs(3293);
    layer1_outputs(3763) <= (layer0_outputs(5859)) and (layer0_outputs(1414));
    layer1_outputs(3764) <= (layer0_outputs(9351)) and not (layer0_outputs(6677));
    layer1_outputs(3765) <= layer0_outputs(8135);
    layer1_outputs(3766) <= not((layer0_outputs(4123)) and (layer0_outputs(4793)));
    layer1_outputs(3767) <= not(layer0_outputs(714)) or (layer0_outputs(1705));
    layer1_outputs(3768) <= '1';
    layer1_outputs(3769) <= not((layer0_outputs(1300)) or (layer0_outputs(1698)));
    layer1_outputs(3770) <= (layer0_outputs(8552)) or (layer0_outputs(3700));
    layer1_outputs(3771) <= not(layer0_outputs(10059));
    layer1_outputs(3772) <= layer0_outputs(3222);
    layer1_outputs(3773) <= not(layer0_outputs(9906)) or (layer0_outputs(8053));
    layer1_outputs(3774) <= layer0_outputs(6069);
    layer1_outputs(3775) <= (layer0_outputs(6741)) and not (layer0_outputs(3315));
    layer1_outputs(3776) <= layer0_outputs(4608);
    layer1_outputs(3777) <= (layer0_outputs(5818)) xor (layer0_outputs(8003));
    layer1_outputs(3778) <= (layer0_outputs(6229)) and not (layer0_outputs(7745));
    layer1_outputs(3779) <= '0';
    layer1_outputs(3780) <= not(layer0_outputs(1869)) or (layer0_outputs(9246));
    layer1_outputs(3781) <= layer0_outputs(9746);
    layer1_outputs(3782) <= layer0_outputs(8763);
    layer1_outputs(3783) <= not(layer0_outputs(8609));
    layer1_outputs(3784) <= (layer0_outputs(3495)) and not (layer0_outputs(1790));
    layer1_outputs(3785) <= (layer0_outputs(2954)) and not (layer0_outputs(9765));
    layer1_outputs(3786) <= not(layer0_outputs(8884)) or (layer0_outputs(9726));
    layer1_outputs(3787) <= (layer0_outputs(3638)) and not (layer0_outputs(5488));
    layer1_outputs(3788) <= not(layer0_outputs(3307));
    layer1_outputs(3789) <= (layer0_outputs(8338)) or (layer0_outputs(3405));
    layer1_outputs(3790) <= (layer0_outputs(6785)) or (layer0_outputs(4745));
    layer1_outputs(3791) <= layer0_outputs(7526);
    layer1_outputs(3792) <= layer0_outputs(657);
    layer1_outputs(3793) <= (layer0_outputs(2026)) and (layer0_outputs(5801));
    layer1_outputs(3794) <= (layer0_outputs(3197)) and not (layer0_outputs(4871));
    layer1_outputs(3795) <= (layer0_outputs(9252)) and not (layer0_outputs(9515));
    layer1_outputs(3796) <= layer0_outputs(2283);
    layer1_outputs(3797) <= not((layer0_outputs(6859)) and (layer0_outputs(9368)));
    layer1_outputs(3798) <= (layer0_outputs(3638)) or (layer0_outputs(7154));
    layer1_outputs(3799) <= not(layer0_outputs(4630)) or (layer0_outputs(1438));
    layer1_outputs(3800) <= layer0_outputs(7512);
    layer1_outputs(3801) <= not(layer0_outputs(5642));
    layer1_outputs(3802) <= layer0_outputs(5049);
    layer1_outputs(3803) <= not((layer0_outputs(538)) and (layer0_outputs(4762)));
    layer1_outputs(3804) <= (layer0_outputs(4981)) and (layer0_outputs(9822));
    layer1_outputs(3805) <= not((layer0_outputs(5467)) or (layer0_outputs(3181)));
    layer1_outputs(3806) <= layer0_outputs(2769);
    layer1_outputs(3807) <= layer0_outputs(2071);
    layer1_outputs(3808) <= (layer0_outputs(3423)) xor (layer0_outputs(4542));
    layer1_outputs(3809) <= (layer0_outputs(1107)) and (layer0_outputs(7864));
    layer1_outputs(3810) <= not(layer0_outputs(9465));
    layer1_outputs(3811) <= layer0_outputs(7441);
    layer1_outputs(3812) <= (layer0_outputs(5327)) and not (layer0_outputs(1015));
    layer1_outputs(3813) <= not((layer0_outputs(2403)) and (layer0_outputs(8283)));
    layer1_outputs(3814) <= not(layer0_outputs(7643)) or (layer0_outputs(6076));
    layer1_outputs(3815) <= '0';
    layer1_outputs(3816) <= not(layer0_outputs(6006));
    layer1_outputs(3817) <= (layer0_outputs(3915)) and not (layer0_outputs(7015));
    layer1_outputs(3818) <= (layer0_outputs(7902)) xor (layer0_outputs(3745));
    layer1_outputs(3819) <= not(layer0_outputs(4196));
    layer1_outputs(3820) <= (layer0_outputs(6064)) xor (layer0_outputs(6520));
    layer1_outputs(3821) <= '1';
    layer1_outputs(3822) <= not((layer0_outputs(6484)) and (layer0_outputs(6681)));
    layer1_outputs(3823) <= (layer0_outputs(9076)) and (layer0_outputs(2394));
    layer1_outputs(3824) <= layer0_outputs(4207);
    layer1_outputs(3825) <= not(layer0_outputs(2899));
    layer1_outputs(3826) <= not((layer0_outputs(5011)) or (layer0_outputs(8086)));
    layer1_outputs(3827) <= (layer0_outputs(5789)) or (layer0_outputs(673));
    layer1_outputs(3828) <= not((layer0_outputs(7849)) and (layer0_outputs(4663)));
    layer1_outputs(3829) <= not(layer0_outputs(7101)) or (layer0_outputs(9520));
    layer1_outputs(3830) <= not((layer0_outputs(7076)) and (layer0_outputs(2076)));
    layer1_outputs(3831) <= not(layer0_outputs(4307)) or (layer0_outputs(412));
    layer1_outputs(3832) <= not(layer0_outputs(8133)) or (layer0_outputs(4084));
    layer1_outputs(3833) <= layer0_outputs(6182);
    layer1_outputs(3834) <= not(layer0_outputs(5179)) or (layer0_outputs(8887));
    layer1_outputs(3835) <= not(layer0_outputs(6450));
    layer1_outputs(3836) <= not(layer0_outputs(4051)) or (layer0_outputs(10073));
    layer1_outputs(3837) <= (layer0_outputs(9000)) or (layer0_outputs(89));
    layer1_outputs(3838) <= (layer0_outputs(9822)) and not (layer0_outputs(9085));
    layer1_outputs(3839) <= not((layer0_outputs(5981)) and (layer0_outputs(3709)));
    layer1_outputs(3840) <= layer0_outputs(6308);
    layer1_outputs(3841) <= (layer0_outputs(7425)) and not (layer0_outputs(9395));
    layer1_outputs(3842) <= not(layer0_outputs(10109)) or (layer0_outputs(6385));
    layer1_outputs(3843) <= '0';
    layer1_outputs(3844) <= '1';
    layer1_outputs(3845) <= not(layer0_outputs(10236));
    layer1_outputs(3846) <= not(layer0_outputs(6428));
    layer1_outputs(3847) <= (layer0_outputs(5863)) and not (layer0_outputs(6497));
    layer1_outputs(3848) <= (layer0_outputs(1921)) and not (layer0_outputs(8339));
    layer1_outputs(3849) <= (layer0_outputs(1497)) or (layer0_outputs(5131));
    layer1_outputs(3850) <= not(layer0_outputs(9921));
    layer1_outputs(3851) <= not((layer0_outputs(7913)) or (layer0_outputs(3750)));
    layer1_outputs(3852) <= (layer0_outputs(454)) and not (layer0_outputs(346));
    layer1_outputs(3853) <= layer0_outputs(3038);
    layer1_outputs(3854) <= not(layer0_outputs(8841)) or (layer0_outputs(1669));
    layer1_outputs(3855) <= (layer0_outputs(411)) and not (layer0_outputs(8738));
    layer1_outputs(3856) <= (layer0_outputs(4462)) and (layer0_outputs(114));
    layer1_outputs(3857) <= layer0_outputs(5181);
    layer1_outputs(3858) <= (layer0_outputs(2652)) or (layer0_outputs(2056));
    layer1_outputs(3859) <= not(layer0_outputs(6266));
    layer1_outputs(3860) <= (layer0_outputs(6186)) and not (layer0_outputs(6393));
    layer1_outputs(3861) <= layer0_outputs(1874);
    layer1_outputs(3862) <= not(layer0_outputs(2509)) or (layer0_outputs(7481));
    layer1_outputs(3863) <= not(layer0_outputs(6139)) or (layer0_outputs(6106));
    layer1_outputs(3864) <= not((layer0_outputs(3914)) and (layer0_outputs(7662)));
    layer1_outputs(3865) <= layer0_outputs(8268);
    layer1_outputs(3866) <= not(layer0_outputs(3393));
    layer1_outputs(3867) <= not((layer0_outputs(3456)) and (layer0_outputs(6283)));
    layer1_outputs(3868) <= not(layer0_outputs(2731));
    layer1_outputs(3869) <= layer0_outputs(5634);
    layer1_outputs(3870) <= (layer0_outputs(8473)) or (layer0_outputs(1772));
    layer1_outputs(3871) <= layer0_outputs(4583);
    layer1_outputs(3872) <= not(layer0_outputs(5719)) or (layer0_outputs(3213));
    layer1_outputs(3873) <= (layer0_outputs(8063)) and not (layer0_outputs(7104));
    layer1_outputs(3874) <= layer0_outputs(4208);
    layer1_outputs(3875) <= not((layer0_outputs(6515)) or (layer0_outputs(3123)));
    layer1_outputs(3876) <= layer0_outputs(4453);
    layer1_outputs(3877) <= layer0_outputs(4284);
    layer1_outputs(3878) <= layer0_outputs(8429);
    layer1_outputs(3879) <= not(layer0_outputs(10117)) or (layer0_outputs(2451));
    layer1_outputs(3880) <= not(layer0_outputs(2473)) or (layer0_outputs(3142));
    layer1_outputs(3881) <= (layer0_outputs(8177)) and not (layer0_outputs(4298));
    layer1_outputs(3882) <= not(layer0_outputs(8215)) or (layer0_outputs(3143));
    layer1_outputs(3883) <= not((layer0_outputs(634)) or (layer0_outputs(9855)));
    layer1_outputs(3884) <= not(layer0_outputs(8838)) or (layer0_outputs(3289));
    layer1_outputs(3885) <= layer0_outputs(2838);
    layer1_outputs(3886) <= not(layer0_outputs(8445));
    layer1_outputs(3887) <= not((layer0_outputs(9566)) or (layer0_outputs(1925)));
    layer1_outputs(3888) <= (layer0_outputs(846)) or (layer0_outputs(9360));
    layer1_outputs(3889) <= not(layer0_outputs(3598)) or (layer0_outputs(7447));
    layer1_outputs(3890) <= (layer0_outputs(6833)) and not (layer0_outputs(7372));
    layer1_outputs(3891) <= '0';
    layer1_outputs(3892) <= '1';
    layer1_outputs(3893) <= (layer0_outputs(6792)) and (layer0_outputs(8665));
    layer1_outputs(3894) <= (layer0_outputs(9910)) and (layer0_outputs(361));
    layer1_outputs(3895) <= layer0_outputs(4576);
    layer1_outputs(3896) <= not(layer0_outputs(5319));
    layer1_outputs(3897) <= not(layer0_outputs(1826));
    layer1_outputs(3898) <= layer0_outputs(1239);
    layer1_outputs(3899) <= layer0_outputs(4280);
    layer1_outputs(3900) <= (layer0_outputs(1230)) and (layer0_outputs(464));
    layer1_outputs(3901) <= '0';
    layer1_outputs(3902) <= not(layer0_outputs(6798)) or (layer0_outputs(8627));
    layer1_outputs(3903) <= layer0_outputs(5815);
    layer1_outputs(3904) <= not(layer0_outputs(8086));
    layer1_outputs(3905) <= not(layer0_outputs(2506)) or (layer0_outputs(3643));
    layer1_outputs(3906) <= '0';
    layer1_outputs(3907) <= not(layer0_outputs(8461));
    layer1_outputs(3908) <= not((layer0_outputs(9729)) and (layer0_outputs(9536)));
    layer1_outputs(3909) <= layer0_outputs(2650);
    layer1_outputs(3910) <= (layer0_outputs(5999)) and (layer0_outputs(2339));
    layer1_outputs(3911) <= (layer0_outputs(753)) and (layer0_outputs(9020));
    layer1_outputs(3912) <= not((layer0_outputs(2062)) or (layer0_outputs(6395)));
    layer1_outputs(3913) <= layer0_outputs(9359);
    layer1_outputs(3914) <= (layer0_outputs(10142)) or (layer0_outputs(9207));
    layer1_outputs(3915) <= not((layer0_outputs(9964)) and (layer0_outputs(9485)));
    layer1_outputs(3916) <= layer0_outputs(2335);
    layer1_outputs(3917) <= not(layer0_outputs(7144)) or (layer0_outputs(3833));
    layer1_outputs(3918) <= layer0_outputs(5201);
    layer1_outputs(3919) <= layer0_outputs(5115);
    layer1_outputs(3920) <= not(layer0_outputs(1262));
    layer1_outputs(3921) <= not(layer0_outputs(7822));
    layer1_outputs(3922) <= layer0_outputs(5046);
    layer1_outputs(3923) <= (layer0_outputs(8734)) and not (layer0_outputs(5387));
    layer1_outputs(3924) <= not((layer0_outputs(2885)) xor (layer0_outputs(1776)));
    layer1_outputs(3925) <= not(layer0_outputs(62)) or (layer0_outputs(3771));
    layer1_outputs(3926) <= not(layer0_outputs(4338)) or (layer0_outputs(7210));
    layer1_outputs(3927) <= (layer0_outputs(3872)) or (layer0_outputs(9012));
    layer1_outputs(3928) <= layer0_outputs(2994);
    layer1_outputs(3929) <= not(layer0_outputs(4351));
    layer1_outputs(3930) <= not(layer0_outputs(10072));
    layer1_outputs(3931) <= (layer0_outputs(6347)) or (layer0_outputs(7549));
    layer1_outputs(3932) <= not(layer0_outputs(1560)) or (layer0_outputs(437));
    layer1_outputs(3933) <= not(layer0_outputs(4684)) or (layer0_outputs(6553));
    layer1_outputs(3934) <= not((layer0_outputs(667)) and (layer0_outputs(489)));
    layer1_outputs(3935) <= not(layer0_outputs(1177)) or (layer0_outputs(1292));
    layer1_outputs(3936) <= (layer0_outputs(6818)) and not (layer0_outputs(517));
    layer1_outputs(3937) <= not(layer0_outputs(5145));
    layer1_outputs(3938) <= (layer0_outputs(4376)) or (layer0_outputs(6368));
    layer1_outputs(3939) <= (layer0_outputs(6388)) or (layer0_outputs(5762));
    layer1_outputs(3940) <= '1';
    layer1_outputs(3941) <= layer0_outputs(419);
    layer1_outputs(3942) <= (layer0_outputs(759)) and (layer0_outputs(8346));
    layer1_outputs(3943) <= layer0_outputs(885);
    layer1_outputs(3944) <= (layer0_outputs(9160)) and not (layer0_outputs(4273));
    layer1_outputs(3945) <= not((layer0_outputs(2828)) and (layer0_outputs(956)));
    layer1_outputs(3946) <= not((layer0_outputs(8007)) xor (layer0_outputs(6312)));
    layer1_outputs(3947) <= (layer0_outputs(7657)) xor (layer0_outputs(8616));
    layer1_outputs(3948) <= not(layer0_outputs(7418)) or (layer0_outputs(5935));
    layer1_outputs(3949) <= not(layer0_outputs(2050)) or (layer0_outputs(5943));
    layer1_outputs(3950) <= '0';
    layer1_outputs(3951) <= (layer0_outputs(8217)) xor (layer0_outputs(1803));
    layer1_outputs(3952) <= '0';
    layer1_outputs(3953) <= not(layer0_outputs(9823));
    layer1_outputs(3954) <= (layer0_outputs(9885)) and not (layer0_outputs(4374));
    layer1_outputs(3955) <= not(layer0_outputs(9839));
    layer1_outputs(3956) <= (layer0_outputs(8651)) and not (layer0_outputs(7527));
    layer1_outputs(3957) <= not((layer0_outputs(1692)) xor (layer0_outputs(2425)));
    layer1_outputs(3958) <= not(layer0_outputs(3610));
    layer1_outputs(3959) <= layer0_outputs(154);
    layer1_outputs(3960) <= (layer0_outputs(2594)) and not (layer0_outputs(2233));
    layer1_outputs(3961) <= not(layer0_outputs(2098)) or (layer0_outputs(3631));
    layer1_outputs(3962) <= (layer0_outputs(4492)) and not (layer0_outputs(1510));
    layer1_outputs(3963) <= not((layer0_outputs(8266)) and (layer0_outputs(7188)));
    layer1_outputs(3964) <= (layer0_outputs(9560)) xor (layer0_outputs(10055));
    layer1_outputs(3965) <= not(layer0_outputs(9354)) or (layer0_outputs(2991));
    layer1_outputs(3966) <= not(layer0_outputs(450));
    layer1_outputs(3967) <= not(layer0_outputs(2893)) or (layer0_outputs(7560));
    layer1_outputs(3968) <= not((layer0_outputs(1060)) and (layer0_outputs(6593)));
    layer1_outputs(3969) <= layer0_outputs(3655);
    layer1_outputs(3970) <= (layer0_outputs(7925)) xor (layer0_outputs(2194));
    layer1_outputs(3971) <= (layer0_outputs(992)) and not (layer0_outputs(2522));
    layer1_outputs(3972) <= not((layer0_outputs(6721)) xor (layer0_outputs(3285)));
    layer1_outputs(3973) <= (layer0_outputs(8973)) and not (layer0_outputs(3407));
    layer1_outputs(3974) <= not((layer0_outputs(5704)) xor (layer0_outputs(9698)));
    layer1_outputs(3975) <= (layer0_outputs(10011)) and not (layer0_outputs(3416));
    layer1_outputs(3976) <= not(layer0_outputs(854));
    layer1_outputs(3977) <= (layer0_outputs(3027)) xor (layer0_outputs(1926));
    layer1_outputs(3978) <= not(layer0_outputs(1636)) or (layer0_outputs(7036));
    layer1_outputs(3979) <= not(layer0_outputs(2492));
    layer1_outputs(3980) <= not(layer0_outputs(3379)) or (layer0_outputs(2757));
    layer1_outputs(3981) <= (layer0_outputs(5088)) and not (layer0_outputs(9648));
    layer1_outputs(3982) <= (layer0_outputs(2730)) xor (layer0_outputs(9014));
    layer1_outputs(3983) <= layer0_outputs(9081);
    layer1_outputs(3984) <= not((layer0_outputs(7076)) and (layer0_outputs(6502)));
    layer1_outputs(3985) <= '1';
    layer1_outputs(3986) <= layer0_outputs(9897);
    layer1_outputs(3987) <= not(layer0_outputs(7658));
    layer1_outputs(3988) <= not((layer0_outputs(6196)) and (layer0_outputs(6418)));
    layer1_outputs(3989) <= layer0_outputs(5943);
    layer1_outputs(3990) <= (layer0_outputs(2809)) and not (layer0_outputs(7704));
    layer1_outputs(3991) <= not(layer0_outputs(10180)) or (layer0_outputs(10052));
    layer1_outputs(3992) <= not(layer0_outputs(3177)) or (layer0_outputs(4710));
    layer1_outputs(3993) <= (layer0_outputs(2153)) and not (layer0_outputs(5483));
    layer1_outputs(3994) <= not((layer0_outputs(1620)) and (layer0_outputs(9345)));
    layer1_outputs(3995) <= not((layer0_outputs(3864)) or (layer0_outputs(3385)));
    layer1_outputs(3996) <= not(layer0_outputs(689));
    layer1_outputs(3997) <= layer0_outputs(5598);
    layer1_outputs(3998) <= not(layer0_outputs(7254));
    layer1_outputs(3999) <= layer0_outputs(6817);
    layer1_outputs(4000) <= (layer0_outputs(6255)) or (layer0_outputs(5023));
    layer1_outputs(4001) <= layer0_outputs(495);
    layer1_outputs(4002) <= (layer0_outputs(5878)) or (layer0_outputs(6746));
    layer1_outputs(4003) <= not(layer0_outputs(2658));
    layer1_outputs(4004) <= not(layer0_outputs(9086));
    layer1_outputs(4005) <= not(layer0_outputs(3283)) or (layer0_outputs(8924));
    layer1_outputs(4006) <= layer0_outputs(1369);
    layer1_outputs(4007) <= (layer0_outputs(3661)) and not (layer0_outputs(9213));
    layer1_outputs(4008) <= not(layer0_outputs(5985));
    layer1_outputs(4009) <= (layer0_outputs(9436)) and not (layer0_outputs(8051));
    layer1_outputs(4010) <= not(layer0_outputs(10127));
    layer1_outputs(4011) <= not((layer0_outputs(1806)) or (layer0_outputs(436)));
    layer1_outputs(4012) <= '1';
    layer1_outputs(4013) <= (layer0_outputs(4167)) and (layer0_outputs(8762));
    layer1_outputs(4014) <= not(layer0_outputs(6082));
    layer1_outputs(4015) <= not((layer0_outputs(1481)) and (layer0_outputs(1189)));
    layer1_outputs(4016) <= (layer0_outputs(7197)) or (layer0_outputs(5865));
    layer1_outputs(4017) <= not(layer0_outputs(4197));
    layer1_outputs(4018) <= (layer0_outputs(6553)) xor (layer0_outputs(5500));
    layer1_outputs(4019) <= not(layer0_outputs(9374)) or (layer0_outputs(9525));
    layer1_outputs(4020) <= not((layer0_outputs(5365)) and (layer0_outputs(3927)));
    layer1_outputs(4021) <= not((layer0_outputs(3669)) or (layer0_outputs(7634)));
    layer1_outputs(4022) <= not((layer0_outputs(4858)) or (layer0_outputs(4345)));
    layer1_outputs(4023) <= (layer0_outputs(6100)) xor (layer0_outputs(6217));
    layer1_outputs(4024) <= not(layer0_outputs(7070));
    layer1_outputs(4025) <= layer0_outputs(8521);
    layer1_outputs(4026) <= not(layer0_outputs(9808));
    layer1_outputs(4027) <= not(layer0_outputs(2719));
    layer1_outputs(4028) <= (layer0_outputs(7797)) and not (layer0_outputs(1827));
    layer1_outputs(4029) <= not(layer0_outputs(6166));
    layer1_outputs(4030) <= not((layer0_outputs(5183)) and (layer0_outputs(6856)));
    layer1_outputs(4031) <= not((layer0_outputs(9673)) or (layer0_outputs(4909)));
    layer1_outputs(4032) <= not((layer0_outputs(1204)) or (layer0_outputs(3449)));
    layer1_outputs(4033) <= layer0_outputs(7928);
    layer1_outputs(4034) <= layer0_outputs(2015);
    layer1_outputs(4035) <= (layer0_outputs(915)) and (layer0_outputs(7224));
    layer1_outputs(4036) <= not((layer0_outputs(3739)) or (layer0_outputs(8284)));
    layer1_outputs(4037) <= not(layer0_outputs(9749));
    layer1_outputs(4038) <= '0';
    layer1_outputs(4039) <= (layer0_outputs(3791)) and not (layer0_outputs(446));
    layer1_outputs(4040) <= not(layer0_outputs(2690));
    layer1_outputs(4041) <= not((layer0_outputs(3330)) and (layer0_outputs(4703)));
    layer1_outputs(4042) <= layer0_outputs(55);
    layer1_outputs(4043) <= (layer0_outputs(342)) and not (layer0_outputs(5053));
    layer1_outputs(4044) <= not((layer0_outputs(9575)) xor (layer0_outputs(7129)));
    layer1_outputs(4045) <= '0';
    layer1_outputs(4046) <= not(layer0_outputs(8397));
    layer1_outputs(4047) <= (layer0_outputs(8634)) or (layer0_outputs(190));
    layer1_outputs(4048) <= layer0_outputs(5562);
    layer1_outputs(4049) <= (layer0_outputs(5271)) or (layer0_outputs(1214));
    layer1_outputs(4050) <= layer0_outputs(1525);
    layer1_outputs(4051) <= not(layer0_outputs(4098)) or (layer0_outputs(6618));
    layer1_outputs(4052) <= layer0_outputs(9887);
    layer1_outputs(4053) <= (layer0_outputs(9637)) or (layer0_outputs(6929));
    layer1_outputs(4054) <= (layer0_outputs(912)) and not (layer0_outputs(7896));
    layer1_outputs(4055) <= (layer0_outputs(6997)) or (layer0_outputs(1562));
    layer1_outputs(4056) <= (layer0_outputs(504)) and not (layer0_outputs(4726));
    layer1_outputs(4057) <= layer0_outputs(8330);
    layer1_outputs(4058) <= not(layer0_outputs(6864));
    layer1_outputs(4059) <= not(layer0_outputs(7798));
    layer1_outputs(4060) <= not(layer0_outputs(1228));
    layer1_outputs(4061) <= not((layer0_outputs(2397)) or (layer0_outputs(2213)));
    layer1_outputs(4062) <= not(layer0_outputs(8614)) or (layer0_outputs(9478));
    layer1_outputs(4063) <= not(layer0_outputs(10115));
    layer1_outputs(4064) <= not((layer0_outputs(153)) or (layer0_outputs(2884)));
    layer1_outputs(4065) <= not(layer0_outputs(9004));
    layer1_outputs(4066) <= not(layer0_outputs(10004));
    layer1_outputs(4067) <= not(layer0_outputs(6313));
    layer1_outputs(4068) <= (layer0_outputs(3846)) or (layer0_outputs(7479));
    layer1_outputs(4069) <= (layer0_outputs(9116)) or (layer0_outputs(1114));
    layer1_outputs(4070) <= not((layer0_outputs(1213)) or (layer0_outputs(467)));
    layer1_outputs(4071) <= not(layer0_outputs(1261));
    layer1_outputs(4072) <= not(layer0_outputs(4254)) or (layer0_outputs(9470));
    layer1_outputs(4073) <= (layer0_outputs(8270)) or (layer0_outputs(1913));
    layer1_outputs(4074) <= not((layer0_outputs(2879)) xor (layer0_outputs(4851)));
    layer1_outputs(4075) <= not((layer0_outputs(6389)) and (layer0_outputs(1721)));
    layer1_outputs(4076) <= layer0_outputs(485);
    layer1_outputs(4077) <= (layer0_outputs(2300)) and not (layer0_outputs(5191));
    layer1_outputs(4078) <= (layer0_outputs(7946)) or (layer0_outputs(1178));
    layer1_outputs(4079) <= layer0_outputs(7179);
    layer1_outputs(4080) <= not(layer0_outputs(1846));
    layer1_outputs(4081) <= not(layer0_outputs(3832)) or (layer0_outputs(10159));
    layer1_outputs(4082) <= not(layer0_outputs(10122)) or (layer0_outputs(3964));
    layer1_outputs(4083) <= (layer0_outputs(6776)) and (layer0_outputs(1506));
    layer1_outputs(4084) <= (layer0_outputs(6022)) xor (layer0_outputs(5268));
    layer1_outputs(4085) <= not(layer0_outputs(8515));
    layer1_outputs(4086) <= not((layer0_outputs(790)) xor (layer0_outputs(1153)));
    layer1_outputs(4087) <= not(layer0_outputs(7962));
    layer1_outputs(4088) <= layer0_outputs(1516);
    layer1_outputs(4089) <= (layer0_outputs(3623)) and not (layer0_outputs(8171));
    layer1_outputs(4090) <= not(layer0_outputs(8367));
    layer1_outputs(4091) <= layer0_outputs(8772);
    layer1_outputs(4092) <= layer0_outputs(9618);
    layer1_outputs(4093) <= not(layer0_outputs(1880)) or (layer0_outputs(794));
    layer1_outputs(4094) <= '0';
    layer1_outputs(4095) <= layer0_outputs(8816);
    layer1_outputs(4096) <= not(layer0_outputs(1536)) or (layer0_outputs(5393));
    layer1_outputs(4097) <= not(layer0_outputs(77));
    layer1_outputs(4098) <= layer0_outputs(7977);
    layer1_outputs(4099) <= (layer0_outputs(9323)) or (layer0_outputs(3730));
    layer1_outputs(4100) <= not((layer0_outputs(7947)) or (layer0_outputs(9490)));
    layer1_outputs(4101) <= layer0_outputs(2460);
    layer1_outputs(4102) <= (layer0_outputs(4151)) and not (layer0_outputs(9701));
    layer1_outputs(4103) <= not(layer0_outputs(8589));
    layer1_outputs(4104) <= not((layer0_outputs(1801)) and (layer0_outputs(7143)));
    layer1_outputs(4105) <= layer0_outputs(1097);
    layer1_outputs(4106) <= (layer0_outputs(2812)) and not (layer0_outputs(4064));
    layer1_outputs(4107) <= not(layer0_outputs(1956)) or (layer0_outputs(5956));
    layer1_outputs(4108) <= not(layer0_outputs(3150));
    layer1_outputs(4109) <= not(layer0_outputs(5307)) or (layer0_outputs(7688));
    layer1_outputs(4110) <= (layer0_outputs(8151)) or (layer0_outputs(4163));
    layer1_outputs(4111) <= not(layer0_outputs(8295));
    layer1_outputs(4112) <= not(layer0_outputs(5889));
    layer1_outputs(4113) <= (layer0_outputs(5968)) xor (layer0_outputs(5668));
    layer1_outputs(4114) <= layer0_outputs(9770);
    layer1_outputs(4115) <= (layer0_outputs(5302)) and (layer0_outputs(1322));
    layer1_outputs(4116) <= not((layer0_outputs(6097)) or (layer0_outputs(2950)));
    layer1_outputs(4117) <= not((layer0_outputs(2806)) and (layer0_outputs(4269)));
    layer1_outputs(4118) <= not(layer0_outputs(3828)) or (layer0_outputs(3221));
    layer1_outputs(4119) <= not(layer0_outputs(6138)) or (layer0_outputs(630));
    layer1_outputs(4120) <= not((layer0_outputs(6473)) or (layer0_outputs(4229)));
    layer1_outputs(4121) <= not(layer0_outputs(8290)) or (layer0_outputs(4305));
    layer1_outputs(4122) <= layer0_outputs(8607);
    layer1_outputs(4123) <= (layer0_outputs(2082)) and not (layer0_outputs(10101));
    layer1_outputs(4124) <= not(layer0_outputs(9981));
    layer1_outputs(4125) <= not((layer0_outputs(9469)) and (layer0_outputs(3860)));
    layer1_outputs(4126) <= (layer0_outputs(2992)) and (layer0_outputs(8283));
    layer1_outputs(4127) <= (layer0_outputs(5363)) and (layer0_outputs(979));
    layer1_outputs(4128) <= not(layer0_outputs(8229));
    layer1_outputs(4129) <= (layer0_outputs(704)) and (layer0_outputs(10079));
    layer1_outputs(4130) <= not(layer0_outputs(9038)) or (layer0_outputs(8810));
    layer1_outputs(4131) <= layer0_outputs(7090);
    layer1_outputs(4132) <= (layer0_outputs(2351)) or (layer0_outputs(488));
    layer1_outputs(4133) <= not(layer0_outputs(1618)) or (layer0_outputs(7301));
    layer1_outputs(4134) <= layer0_outputs(4721);
    layer1_outputs(4135) <= not((layer0_outputs(8647)) xor (layer0_outputs(3173)));
    layer1_outputs(4136) <= layer0_outputs(2613);
    layer1_outputs(4137) <= layer0_outputs(6536);
    layer1_outputs(4138) <= layer0_outputs(4962);
    layer1_outputs(4139) <= not(layer0_outputs(8963));
    layer1_outputs(4140) <= not(layer0_outputs(4040));
    layer1_outputs(4141) <= not(layer0_outputs(2937));
    layer1_outputs(4142) <= '1';
    layer1_outputs(4143) <= '0';
    layer1_outputs(4144) <= not(layer0_outputs(6093));
    layer1_outputs(4145) <= (layer0_outputs(822)) and not (layer0_outputs(397));
    layer1_outputs(4146) <= layer0_outputs(827);
    layer1_outputs(4147) <= (layer0_outputs(6757)) or (layer0_outputs(2656));
    layer1_outputs(4148) <= (layer0_outputs(10208)) and not (layer0_outputs(2332));
    layer1_outputs(4149) <= not(layer0_outputs(2497)) or (layer0_outputs(750));
    layer1_outputs(4150) <= (layer0_outputs(5509)) and not (layer0_outputs(3025));
    layer1_outputs(4151) <= not((layer0_outputs(4065)) or (layer0_outputs(9577)));
    layer1_outputs(4152) <= not(layer0_outputs(3978)) or (layer0_outputs(1428));
    layer1_outputs(4153) <= not((layer0_outputs(6655)) and (layer0_outputs(1724)));
    layer1_outputs(4154) <= not((layer0_outputs(1162)) or (layer0_outputs(2561)));
    layer1_outputs(4155) <= not(layer0_outputs(4845)) or (layer0_outputs(9725));
    layer1_outputs(4156) <= layer0_outputs(4429);
    layer1_outputs(4157) <= (layer0_outputs(7668)) and not (layer0_outputs(371));
    layer1_outputs(4158) <= layer0_outputs(1351);
    layer1_outputs(4159) <= not(layer0_outputs(7737));
    layer1_outputs(4160) <= not((layer0_outputs(119)) and (layer0_outputs(9313)));
    layer1_outputs(4161) <= layer0_outputs(717);
    layer1_outputs(4162) <= not((layer0_outputs(7587)) and (layer0_outputs(8478)));
    layer1_outputs(4163) <= layer0_outputs(9874);
    layer1_outputs(4164) <= not(layer0_outputs(1796)) or (layer0_outputs(9439));
    layer1_outputs(4165) <= not(layer0_outputs(6501));
    layer1_outputs(4166) <= not(layer0_outputs(5076));
    layer1_outputs(4167) <= not(layer0_outputs(3916));
    layer1_outputs(4168) <= layer0_outputs(7657);
    layer1_outputs(4169) <= not(layer0_outputs(7887));
    layer1_outputs(4170) <= (layer0_outputs(271)) and (layer0_outputs(1351));
    layer1_outputs(4171) <= (layer0_outputs(4020)) and (layer0_outputs(1676));
    layer1_outputs(4172) <= layer0_outputs(210);
    layer1_outputs(4173) <= (layer0_outputs(2388)) or (layer0_outputs(10209));
    layer1_outputs(4174) <= not((layer0_outputs(6349)) or (layer0_outputs(8398)));
    layer1_outputs(4175) <= not((layer0_outputs(6826)) or (layer0_outputs(5216)));
    layer1_outputs(4176) <= not((layer0_outputs(3196)) xor (layer0_outputs(2537)));
    layer1_outputs(4177) <= (layer0_outputs(8306)) and not (layer0_outputs(5426));
    layer1_outputs(4178) <= not(layer0_outputs(7008)) or (layer0_outputs(3895));
    layer1_outputs(4179) <= not((layer0_outputs(346)) xor (layer0_outputs(534)));
    layer1_outputs(4180) <= not(layer0_outputs(4032));
    layer1_outputs(4181) <= layer0_outputs(1875);
    layer1_outputs(4182) <= not((layer0_outputs(4103)) and (layer0_outputs(9853)));
    layer1_outputs(4183) <= not(layer0_outputs(1416)) or (layer0_outputs(3043));
    layer1_outputs(4184) <= '0';
    layer1_outputs(4185) <= (layer0_outputs(10076)) or (layer0_outputs(3097));
    layer1_outputs(4186) <= not(layer0_outputs(4785)) or (layer0_outputs(1336));
    layer1_outputs(4187) <= layer0_outputs(806);
    layer1_outputs(4188) <= (layer0_outputs(7147)) and not (layer0_outputs(6630));
    layer1_outputs(4189) <= (layer0_outputs(8018)) xor (layer0_outputs(4336));
    layer1_outputs(4190) <= not(layer0_outputs(10013));
    layer1_outputs(4191) <= layer0_outputs(4490);
    layer1_outputs(4192) <= layer0_outputs(10175);
    layer1_outputs(4193) <= layer0_outputs(6373);
    layer1_outputs(4194) <= (layer0_outputs(7606)) and not (layer0_outputs(1665));
    layer1_outputs(4195) <= not(layer0_outputs(2048));
    layer1_outputs(4196) <= not(layer0_outputs(1226));
    layer1_outputs(4197) <= (layer0_outputs(4318)) and not (layer0_outputs(3374));
    layer1_outputs(4198) <= not(layer0_outputs(3091));
    layer1_outputs(4199) <= (layer0_outputs(1427)) and not (layer0_outputs(1341));
    layer1_outputs(4200) <= not((layer0_outputs(5415)) or (layer0_outputs(9886)));
    layer1_outputs(4201) <= not((layer0_outputs(2192)) and (layer0_outputs(8221)));
    layer1_outputs(4202) <= (layer0_outputs(1895)) xor (layer0_outputs(749));
    layer1_outputs(4203) <= layer0_outputs(3754);
    layer1_outputs(4204) <= layer0_outputs(550);
    layer1_outputs(4205) <= not(layer0_outputs(5006)) or (layer0_outputs(985));
    layer1_outputs(4206) <= (layer0_outputs(6888)) xor (layer0_outputs(6229));
    layer1_outputs(4207) <= layer0_outputs(4772);
    layer1_outputs(4208) <= not((layer0_outputs(5769)) xor (layer0_outputs(10056)));
    layer1_outputs(4209) <= layer0_outputs(410);
    layer1_outputs(4210) <= not((layer0_outputs(7435)) xor (layer0_outputs(904)));
    layer1_outputs(4211) <= (layer0_outputs(3508)) and (layer0_outputs(2655));
    layer1_outputs(4212) <= not((layer0_outputs(4775)) or (layer0_outputs(7944)));
    layer1_outputs(4213) <= not(layer0_outputs(4872));
    layer1_outputs(4214) <= (layer0_outputs(5510)) and not (layer0_outputs(1986));
    layer1_outputs(4215) <= (layer0_outputs(7920)) or (layer0_outputs(6532));
    layer1_outputs(4216) <= not(layer0_outputs(4906)) or (layer0_outputs(4062));
    layer1_outputs(4217) <= not(layer0_outputs(4976));
    layer1_outputs(4218) <= not(layer0_outputs(7222)) or (layer0_outputs(8430));
    layer1_outputs(4219) <= layer0_outputs(2928);
    layer1_outputs(4220) <= not((layer0_outputs(7159)) or (layer0_outputs(7971)));
    layer1_outputs(4221) <= not(layer0_outputs(8861)) or (layer0_outputs(2065));
    layer1_outputs(4222) <= '0';
    layer1_outputs(4223) <= not(layer0_outputs(3296));
    layer1_outputs(4224) <= not((layer0_outputs(6882)) xor (layer0_outputs(5371)));
    layer1_outputs(4225) <= layer0_outputs(8988);
    layer1_outputs(4226) <= (layer0_outputs(2067)) and not (layer0_outputs(10007));
    layer1_outputs(4227) <= not(layer0_outputs(120));
    layer1_outputs(4228) <= layer0_outputs(2211);
    layer1_outputs(4229) <= (layer0_outputs(2886)) and (layer0_outputs(5075));
    layer1_outputs(4230) <= not((layer0_outputs(3248)) or (layer0_outputs(830)));
    layer1_outputs(4231) <= not(layer0_outputs(2208));
    layer1_outputs(4232) <= not(layer0_outputs(5121));
    layer1_outputs(4233) <= not(layer0_outputs(3534));
    layer1_outputs(4234) <= not(layer0_outputs(9979));
    layer1_outputs(4235) <= layer0_outputs(2520);
    layer1_outputs(4236) <= (layer0_outputs(1438)) and not (layer0_outputs(9997));
    layer1_outputs(4237) <= (layer0_outputs(6752)) or (layer0_outputs(5869));
    layer1_outputs(4238) <= not((layer0_outputs(2953)) or (layer0_outputs(7217)));
    layer1_outputs(4239) <= not(layer0_outputs(244));
    layer1_outputs(4240) <= layer0_outputs(4460);
    layer1_outputs(4241) <= layer0_outputs(5886);
    layer1_outputs(4242) <= not((layer0_outputs(1466)) or (layer0_outputs(1808)));
    layer1_outputs(4243) <= not(layer0_outputs(4831)) or (layer0_outputs(7459));
    layer1_outputs(4244) <= not(layer0_outputs(5269)) or (layer0_outputs(41));
    layer1_outputs(4245) <= (layer0_outputs(8269)) and not (layer0_outputs(8202));
    layer1_outputs(4246) <= layer0_outputs(3016);
    layer1_outputs(4247) <= not((layer0_outputs(7516)) and (layer0_outputs(2262)));
    layer1_outputs(4248) <= layer0_outputs(10155);
    layer1_outputs(4249) <= layer0_outputs(2116);
    layer1_outputs(4250) <= not(layer0_outputs(8276)) or (layer0_outputs(1999));
    layer1_outputs(4251) <= layer0_outputs(4517);
    layer1_outputs(4252) <= not((layer0_outputs(5379)) or (layer0_outputs(475)));
    layer1_outputs(4253) <= layer0_outputs(5988);
    layer1_outputs(4254) <= (layer0_outputs(334)) and not (layer0_outputs(3888));
    layer1_outputs(4255) <= layer0_outputs(405);
    layer1_outputs(4256) <= (layer0_outputs(4215)) and (layer0_outputs(10019));
    layer1_outputs(4257) <= (layer0_outputs(5134)) and not (layer0_outputs(3105));
    layer1_outputs(4258) <= not(layer0_outputs(7975));
    layer1_outputs(4259) <= not(layer0_outputs(7984));
    layer1_outputs(4260) <= not(layer0_outputs(1144)) or (layer0_outputs(6243));
    layer1_outputs(4261) <= (layer0_outputs(1211)) and not (layer0_outputs(1401));
    layer1_outputs(4262) <= not(layer0_outputs(5108));
    layer1_outputs(4263) <= not(layer0_outputs(411));
    layer1_outputs(4264) <= layer0_outputs(8094);
    layer1_outputs(4265) <= (layer0_outputs(540)) and (layer0_outputs(7007));
    layer1_outputs(4266) <= not(layer0_outputs(5135));
    layer1_outputs(4267) <= not((layer0_outputs(1679)) xor (layer0_outputs(1753)));
    layer1_outputs(4268) <= not(layer0_outputs(679)) or (layer0_outputs(6472));
    layer1_outputs(4269) <= not(layer0_outputs(1188));
    layer1_outputs(4270) <= (layer0_outputs(9517)) and not (layer0_outputs(3107));
    layer1_outputs(4271) <= not(layer0_outputs(4180));
    layer1_outputs(4272) <= not(layer0_outputs(9883));
    layer1_outputs(4273) <= (layer0_outputs(6773)) and (layer0_outputs(1360));
    layer1_outputs(4274) <= '1';
    layer1_outputs(4275) <= (layer0_outputs(9652)) and not (layer0_outputs(4380));
    layer1_outputs(4276) <= layer0_outputs(4378);
    layer1_outputs(4277) <= (layer0_outputs(7627)) xor (layer0_outputs(3417));
    layer1_outputs(4278) <= (layer0_outputs(1919)) or (layer0_outputs(2906));
    layer1_outputs(4279) <= (layer0_outputs(9569)) and not (layer0_outputs(1577));
    layer1_outputs(4280) <= not(layer0_outputs(5032));
    layer1_outputs(4281) <= layer0_outputs(3863);
    layer1_outputs(4282) <= layer0_outputs(4771);
    layer1_outputs(4283) <= not(layer0_outputs(3330));
    layer1_outputs(4284) <= (layer0_outputs(5950)) or (layer0_outputs(8990));
    layer1_outputs(4285) <= (layer0_outputs(878)) or (layer0_outputs(4914));
    layer1_outputs(4286) <= not(layer0_outputs(5888)) or (layer0_outputs(4589));
    layer1_outputs(4287) <= layer0_outputs(9866);
    layer1_outputs(4288) <= (layer0_outputs(7707)) xor (layer0_outputs(3966));
    layer1_outputs(4289) <= not(layer0_outputs(305)) or (layer0_outputs(5790));
    layer1_outputs(4290) <= not(layer0_outputs(7078));
    layer1_outputs(4291) <= (layer0_outputs(5062)) and (layer0_outputs(1712));
    layer1_outputs(4292) <= layer0_outputs(2289);
    layer1_outputs(4293) <= layer0_outputs(3334);
    layer1_outputs(4294) <= layer0_outputs(6498);
    layer1_outputs(4295) <= (layer0_outputs(5469)) and not (layer0_outputs(4949));
    layer1_outputs(4296) <= not(layer0_outputs(7392)) or (layer0_outputs(9903));
    layer1_outputs(4297) <= layer0_outputs(4194);
    layer1_outputs(4298) <= (layer0_outputs(5811)) and not (layer0_outputs(921));
    layer1_outputs(4299) <= not((layer0_outputs(4069)) or (layer0_outputs(5843)));
    layer1_outputs(4300) <= not((layer0_outputs(8812)) or (layer0_outputs(9468)));
    layer1_outputs(4301) <= layer0_outputs(8064);
    layer1_outputs(4302) <= (layer0_outputs(1938)) and not (layer0_outputs(5585));
    layer1_outputs(4303) <= not(layer0_outputs(1591));
    layer1_outputs(4304) <= (layer0_outputs(455)) xor (layer0_outputs(3920));
    layer1_outputs(4305) <= not(layer0_outputs(7216));
    layer1_outputs(4306) <= '1';
    layer1_outputs(4307) <= layer0_outputs(5067);
    layer1_outputs(4308) <= (layer0_outputs(8970)) xor (layer0_outputs(596));
    layer1_outputs(4309) <= not(layer0_outputs(5890)) or (layer0_outputs(1511));
    layer1_outputs(4310) <= not(layer0_outputs(4751));
    layer1_outputs(4311) <= (layer0_outputs(9528)) or (layer0_outputs(4537));
    layer1_outputs(4312) <= (layer0_outputs(8300)) and not (layer0_outputs(9723));
    layer1_outputs(4313) <= not(layer0_outputs(1848));
    layer1_outputs(4314) <= layer0_outputs(5236);
    layer1_outputs(4315) <= layer0_outputs(1234);
    layer1_outputs(4316) <= not((layer0_outputs(8181)) or (layer0_outputs(35)));
    layer1_outputs(4317) <= not(layer0_outputs(9178)) or (layer0_outputs(618));
    layer1_outputs(4318) <= not(layer0_outputs(8701)) or (layer0_outputs(7450));
    layer1_outputs(4319) <= not(layer0_outputs(2092));
    layer1_outputs(4320) <= '0';
    layer1_outputs(4321) <= (layer0_outputs(8505)) xor (layer0_outputs(9274));
    layer1_outputs(4322) <= layer0_outputs(1189);
    layer1_outputs(4323) <= (layer0_outputs(3154)) and (layer0_outputs(7387));
    layer1_outputs(4324) <= not((layer0_outputs(6145)) and (layer0_outputs(9235)));
    layer1_outputs(4325) <= (layer0_outputs(3811)) and not (layer0_outputs(8915));
    layer1_outputs(4326) <= (layer0_outputs(3211)) and not (layer0_outputs(7112));
    layer1_outputs(4327) <= layer0_outputs(8079);
    layer1_outputs(4328) <= layer0_outputs(5711);
    layer1_outputs(4329) <= not(layer0_outputs(7398));
    layer1_outputs(4330) <= not(layer0_outputs(4630));
    layer1_outputs(4331) <= not(layer0_outputs(8295));
    layer1_outputs(4332) <= layer0_outputs(6558);
    layer1_outputs(4333) <= (layer0_outputs(3905)) and not (layer0_outputs(1548));
    layer1_outputs(4334) <= (layer0_outputs(989)) xor (layer0_outputs(3919));
    layer1_outputs(4335) <= not((layer0_outputs(8829)) xor (layer0_outputs(8599)));
    layer1_outputs(4336) <= not(layer0_outputs(663));
    layer1_outputs(4337) <= not((layer0_outputs(2144)) xor (layer0_outputs(8405)));
    layer1_outputs(4338) <= not(layer0_outputs(4716));
    layer1_outputs(4339) <= (layer0_outputs(8329)) or (layer0_outputs(4608));
    layer1_outputs(4340) <= not((layer0_outputs(5231)) and (layer0_outputs(935)));
    layer1_outputs(4341) <= not(layer0_outputs(2804)) or (layer0_outputs(2683));
    layer1_outputs(4342) <= not(layer0_outputs(3612));
    layer1_outputs(4343) <= (layer0_outputs(9556)) and (layer0_outputs(3063));
    layer1_outputs(4344) <= not(layer0_outputs(1015));
    layer1_outputs(4345) <= layer0_outputs(9421);
    layer1_outputs(4346) <= (layer0_outputs(5452)) and not (layer0_outputs(2959));
    layer1_outputs(4347) <= '1';
    layer1_outputs(4348) <= layer0_outputs(8345);
    layer1_outputs(4349) <= layer0_outputs(2806);
    layer1_outputs(4350) <= (layer0_outputs(7824)) or (layer0_outputs(294));
    layer1_outputs(4351) <= not((layer0_outputs(9472)) or (layer0_outputs(6471)));
    layer1_outputs(4352) <= layer0_outputs(6968);
    layer1_outputs(4353) <= (layer0_outputs(8315)) and not (layer0_outputs(8978));
    layer1_outputs(4354) <= (layer0_outputs(2996)) and not (layer0_outputs(2478));
    layer1_outputs(4355) <= not((layer0_outputs(3842)) and (layer0_outputs(8317)));
    layer1_outputs(4356) <= not((layer0_outputs(9736)) xor (layer0_outputs(1658)));
    layer1_outputs(4357) <= not((layer0_outputs(7496)) or (layer0_outputs(3006)));
    layer1_outputs(4358) <= (layer0_outputs(104)) or (layer0_outputs(3360));
    layer1_outputs(4359) <= '1';
    layer1_outputs(4360) <= not(layer0_outputs(6219));
    layer1_outputs(4361) <= (layer0_outputs(4025)) or (layer0_outputs(732));
    layer1_outputs(4362) <= (layer0_outputs(8857)) and (layer0_outputs(10216));
    layer1_outputs(4363) <= not((layer0_outputs(1862)) or (layer0_outputs(5856)));
    layer1_outputs(4364) <= not(layer0_outputs(3286)) or (layer0_outputs(4732));
    layer1_outputs(4365) <= not((layer0_outputs(523)) xor (layer0_outputs(8881)));
    layer1_outputs(4366) <= '1';
    layer1_outputs(4367) <= not(layer0_outputs(2802));
    layer1_outputs(4368) <= layer0_outputs(9032);
    layer1_outputs(4369) <= not(layer0_outputs(8374));
    layer1_outputs(4370) <= not((layer0_outputs(6949)) xor (layer0_outputs(3765)));
    layer1_outputs(4371) <= (layer0_outputs(9630)) and (layer0_outputs(2867));
    layer1_outputs(4372) <= not((layer0_outputs(1689)) xor (layer0_outputs(1510)));
    layer1_outputs(4373) <= layer0_outputs(7637);
    layer1_outputs(4374) <= (layer0_outputs(6345)) xor (layer0_outputs(5334));
    layer1_outputs(4375) <= not(layer0_outputs(7611));
    layer1_outputs(4376) <= not(layer0_outputs(4067));
    layer1_outputs(4377) <= layer0_outputs(4894);
    layer1_outputs(4378) <= not((layer0_outputs(8043)) or (layer0_outputs(4884)));
    layer1_outputs(4379) <= '1';
    layer1_outputs(4380) <= (layer0_outputs(4635)) and not (layer0_outputs(5331));
    layer1_outputs(4381) <= not(layer0_outputs(9147));
    layer1_outputs(4382) <= (layer0_outputs(6874)) and (layer0_outputs(7056));
    layer1_outputs(4383) <= layer0_outputs(8092);
    layer1_outputs(4384) <= (layer0_outputs(10042)) xor (layer0_outputs(5838));
    layer1_outputs(4385) <= not(layer0_outputs(6979));
    layer1_outputs(4386) <= (layer0_outputs(6056)) and (layer0_outputs(3546));
    layer1_outputs(4387) <= (layer0_outputs(8443)) and (layer0_outputs(6367));
    layer1_outputs(4388) <= not((layer0_outputs(5072)) or (layer0_outputs(546)));
    layer1_outputs(4389) <= not((layer0_outputs(4323)) and (layer0_outputs(235)));
    layer1_outputs(4390) <= (layer0_outputs(386)) and not (layer0_outputs(2123));
    layer1_outputs(4391) <= (layer0_outputs(8071)) and (layer0_outputs(2727));
    layer1_outputs(4392) <= not((layer0_outputs(1513)) or (layer0_outputs(6791)));
    layer1_outputs(4393) <= layer0_outputs(1283);
    layer1_outputs(4394) <= layer0_outputs(3191);
    layer1_outputs(4395) <= (layer0_outputs(249)) or (layer0_outputs(1375));
    layer1_outputs(4396) <= not(layer0_outputs(5862));
    layer1_outputs(4397) <= not((layer0_outputs(7855)) xor (layer0_outputs(2510)));
    layer1_outputs(4398) <= (layer0_outputs(3725)) or (layer0_outputs(5735));
    layer1_outputs(4399) <= layer0_outputs(6420);
    layer1_outputs(4400) <= not(layer0_outputs(5228)) or (layer0_outputs(9524));
    layer1_outputs(4401) <= not(layer0_outputs(6901)) or (layer0_outputs(5131));
    layer1_outputs(4402) <= not((layer0_outputs(4101)) and (layer0_outputs(9657)));
    layer1_outputs(4403) <= layer0_outputs(7112);
    layer1_outputs(4404) <= not(layer0_outputs(4144)) or (layer0_outputs(10062));
    layer1_outputs(4405) <= not((layer0_outputs(5698)) and (layer0_outputs(8755)));
    layer1_outputs(4406) <= not((layer0_outputs(5405)) and (layer0_outputs(1935)));
    layer1_outputs(4407) <= not(layer0_outputs(736));
    layer1_outputs(4408) <= (layer0_outputs(4674)) and not (layer0_outputs(5612));
    layer1_outputs(4409) <= (layer0_outputs(1470)) xor (layer0_outputs(2960));
    layer1_outputs(4410) <= (layer0_outputs(752)) and not (layer0_outputs(4688));
    layer1_outputs(4411) <= not((layer0_outputs(2148)) and (layer0_outputs(9534)));
    layer1_outputs(4412) <= (layer0_outputs(4893)) and not (layer0_outputs(5567));
    layer1_outputs(4413) <= layer0_outputs(8776);
    layer1_outputs(4414) <= (layer0_outputs(6572)) xor (layer0_outputs(1264));
    layer1_outputs(4415) <= not(layer0_outputs(5262));
    layer1_outputs(4416) <= (layer0_outputs(4205)) and not (layer0_outputs(2321));
    layer1_outputs(4417) <= not((layer0_outputs(6315)) or (layer0_outputs(4802)));
    layer1_outputs(4418) <= layer0_outputs(5516);
    layer1_outputs(4419) <= not(layer0_outputs(3532));
    layer1_outputs(4420) <= not(layer0_outputs(5977));
    layer1_outputs(4421) <= not((layer0_outputs(4521)) and (layer0_outputs(1939)));
    layer1_outputs(4422) <= (layer0_outputs(4468)) and (layer0_outputs(7461));
    layer1_outputs(4423) <= (layer0_outputs(1149)) and not (layer0_outputs(1938));
    layer1_outputs(4424) <= (layer0_outputs(1731)) and (layer0_outputs(1315));
    layer1_outputs(4425) <= not(layer0_outputs(8547)) or (layer0_outputs(6383));
    layer1_outputs(4426) <= not(layer0_outputs(7242));
    layer1_outputs(4427) <= (layer0_outputs(9936)) and not (layer0_outputs(2966));
    layer1_outputs(4428) <= not(layer0_outputs(2038)) or (layer0_outputs(4186));
    layer1_outputs(4429) <= layer0_outputs(3288);
    layer1_outputs(4430) <= not(layer0_outputs(1882));
    layer1_outputs(4431) <= (layer0_outputs(8476)) or (layer0_outputs(9138));
    layer1_outputs(4432) <= not(layer0_outputs(6259));
    layer1_outputs(4433) <= '1';
    layer1_outputs(4434) <= not(layer0_outputs(7977));
    layer1_outputs(4435) <= not(layer0_outputs(9994)) or (layer0_outputs(9846));
    layer1_outputs(4436) <= not(layer0_outputs(541));
    layer1_outputs(4437) <= not(layer0_outputs(5257)) or (layer0_outputs(3264));
    layer1_outputs(4438) <= not(layer0_outputs(5431));
    layer1_outputs(4439) <= not(layer0_outputs(1219));
    layer1_outputs(4440) <= not((layer0_outputs(2072)) xor (layer0_outputs(4243)));
    layer1_outputs(4441) <= not((layer0_outputs(3382)) or (layer0_outputs(5515)));
    layer1_outputs(4442) <= not(layer0_outputs(6645));
    layer1_outputs(4443) <= not((layer0_outputs(3541)) xor (layer0_outputs(957)));
    layer1_outputs(4444) <= layer0_outputs(1803);
    layer1_outputs(4445) <= not((layer0_outputs(964)) xor (layer0_outputs(7278)));
    layer1_outputs(4446) <= not(layer0_outputs(3882));
    layer1_outputs(4447) <= not((layer0_outputs(5102)) xor (layer0_outputs(4699)));
    layer1_outputs(4448) <= '0';
    layer1_outputs(4449) <= not((layer0_outputs(9033)) and (layer0_outputs(2743)));
    layer1_outputs(4450) <= not(layer0_outputs(4567)) or (layer0_outputs(5278));
    layer1_outputs(4451) <= (layer0_outputs(7876)) and (layer0_outputs(7142));
    layer1_outputs(4452) <= (layer0_outputs(3932)) xor (layer0_outputs(1589));
    layer1_outputs(4453) <= layer0_outputs(2527);
    layer1_outputs(4454) <= not(layer0_outputs(6545));
    layer1_outputs(4455) <= (layer0_outputs(3136)) and not (layer0_outputs(16));
    layer1_outputs(4456) <= not(layer0_outputs(9871)) or (layer0_outputs(1268));
    layer1_outputs(4457) <= not((layer0_outputs(465)) or (layer0_outputs(4786)));
    layer1_outputs(4458) <= not((layer0_outputs(10070)) xor (layer0_outputs(8246)));
    layer1_outputs(4459) <= not(layer0_outputs(9069)) or (layer0_outputs(8134));
    layer1_outputs(4460) <= layer0_outputs(997);
    layer1_outputs(4461) <= not((layer0_outputs(6661)) or (layer0_outputs(5625)));
    layer1_outputs(4462) <= (layer0_outputs(7801)) and not (layer0_outputs(2601));
    layer1_outputs(4463) <= not(layer0_outputs(1475)) or (layer0_outputs(9160));
    layer1_outputs(4464) <= not(layer0_outputs(4389));
    layer1_outputs(4465) <= (layer0_outputs(5397)) xor (layer0_outputs(9487));
    layer1_outputs(4466) <= (layer0_outputs(6836)) xor (layer0_outputs(2557));
    layer1_outputs(4467) <= '1';
    layer1_outputs(4468) <= layer0_outputs(6409);
    layer1_outputs(4469) <= (layer0_outputs(8995)) or (layer0_outputs(2729));
    layer1_outputs(4470) <= not(layer0_outputs(4519)) or (layer0_outputs(8542));
    layer1_outputs(4471) <= (layer0_outputs(3433)) xor (layer0_outputs(6293));
    layer1_outputs(4472) <= not(layer0_outputs(5477));
    layer1_outputs(4473) <= not((layer0_outputs(1077)) xor (layer0_outputs(4862)));
    layer1_outputs(4474) <= layer0_outputs(5427);
    layer1_outputs(4475) <= (layer0_outputs(5007)) and not (layer0_outputs(8460));
    layer1_outputs(4476) <= not((layer0_outputs(2105)) or (layer0_outputs(1819)));
    layer1_outputs(4477) <= (layer0_outputs(145)) and not (layer0_outputs(8687));
    layer1_outputs(4478) <= not((layer0_outputs(7769)) and (layer0_outputs(6749)));
    layer1_outputs(4479) <= (layer0_outputs(372)) and not (layer0_outputs(3352));
    layer1_outputs(4480) <= layer0_outputs(9295);
    layer1_outputs(4481) <= not(layer0_outputs(3510)) or (layer0_outputs(3962));
    layer1_outputs(4482) <= not(layer0_outputs(7371)) or (layer0_outputs(10120));
    layer1_outputs(4483) <= not(layer0_outputs(63)) or (layer0_outputs(6422));
    layer1_outputs(4484) <= not(layer0_outputs(417)) or (layer0_outputs(6528));
    layer1_outputs(4485) <= not(layer0_outputs(1359));
    layer1_outputs(4486) <= layer0_outputs(5534);
    layer1_outputs(4487) <= (layer0_outputs(2986)) xor (layer0_outputs(1236));
    layer1_outputs(4488) <= layer0_outputs(2074);
    layer1_outputs(4489) <= '1';
    layer1_outputs(4490) <= (layer0_outputs(8267)) and (layer0_outputs(6966));
    layer1_outputs(4491) <= not(layer0_outputs(2880)) or (layer0_outputs(6571));
    layer1_outputs(4492) <= (layer0_outputs(5361)) or (layer0_outputs(2030));
    layer1_outputs(4493) <= (layer0_outputs(6415)) and (layer0_outputs(9349));
    layer1_outputs(4494) <= not(layer0_outputs(4609)) or (layer0_outputs(4702));
    layer1_outputs(4495) <= not(layer0_outputs(9471)) or (layer0_outputs(5562));
    layer1_outputs(4496) <= (layer0_outputs(6213)) or (layer0_outputs(1749));
    layer1_outputs(4497) <= not(layer0_outputs(9689));
    layer1_outputs(4498) <= not(layer0_outputs(9339));
    layer1_outputs(4499) <= not(layer0_outputs(9516));
    layer1_outputs(4500) <= not(layer0_outputs(4987));
    layer1_outputs(4501) <= not((layer0_outputs(5721)) or (layer0_outputs(9012)));
    layer1_outputs(4502) <= layer0_outputs(1249);
    layer1_outputs(4503) <= not(layer0_outputs(4948));
    layer1_outputs(4504) <= (layer0_outputs(2001)) xor (layer0_outputs(1854));
    layer1_outputs(4505) <= (layer0_outputs(3679)) xor (layer0_outputs(8835));
    layer1_outputs(4506) <= not(layer0_outputs(4212)) or (layer0_outputs(9747));
    layer1_outputs(4507) <= not(layer0_outputs(4454));
    layer1_outputs(4508) <= not(layer0_outputs(6397));
    layer1_outputs(4509) <= not(layer0_outputs(4539)) or (layer0_outputs(629));
    layer1_outputs(4510) <= '1';
    layer1_outputs(4511) <= (layer0_outputs(8632)) or (layer0_outputs(1992));
    layer1_outputs(4512) <= (layer0_outputs(5472)) xor (layer0_outputs(4678));
    layer1_outputs(4513) <= not((layer0_outputs(9544)) or (layer0_outputs(7653)));
    layer1_outputs(4514) <= (layer0_outputs(2284)) or (layer0_outputs(6619));
    layer1_outputs(4515) <= (layer0_outputs(1964)) or (layer0_outputs(7666));
    layer1_outputs(4516) <= layer0_outputs(5119);
    layer1_outputs(4517) <= not(layer0_outputs(10067));
    layer1_outputs(4518) <= layer0_outputs(8977);
    layer1_outputs(4519) <= not(layer0_outputs(4061)) or (layer0_outputs(2967));
    layer1_outputs(4520) <= '1';
    layer1_outputs(4521) <= (layer0_outputs(5739)) xor (layer0_outputs(2758));
    layer1_outputs(4522) <= layer0_outputs(1994);
    layer1_outputs(4523) <= not(layer0_outputs(8957)) or (layer0_outputs(2602));
    layer1_outputs(4524) <= not(layer0_outputs(5913));
    layer1_outputs(4525) <= not(layer0_outputs(9250));
    layer1_outputs(4526) <= (layer0_outputs(4126)) or (layer0_outputs(3483));
    layer1_outputs(4527) <= '1';
    layer1_outputs(4528) <= not((layer0_outputs(5187)) and (layer0_outputs(4416)));
    layer1_outputs(4529) <= not(layer0_outputs(5528));
    layer1_outputs(4530) <= (layer0_outputs(826)) and not (layer0_outputs(685));
    layer1_outputs(4531) <= layer0_outputs(1469);
    layer1_outputs(4532) <= layer0_outputs(7456);
    layer1_outputs(4533) <= not(layer0_outputs(5852)) or (layer0_outputs(4546));
    layer1_outputs(4534) <= layer0_outputs(7573);
    layer1_outputs(4535) <= not((layer0_outputs(4755)) and (layer0_outputs(1652)));
    layer1_outputs(4536) <= not(layer0_outputs(2458)) or (layer0_outputs(1352));
    layer1_outputs(4537) <= (layer0_outputs(7407)) and not (layer0_outputs(7817));
    layer1_outputs(4538) <= not(layer0_outputs(9852)) or (layer0_outputs(9837));
    layer1_outputs(4539) <= layer0_outputs(4187);
    layer1_outputs(4540) <= layer0_outputs(6263);
    layer1_outputs(4541) <= not(layer0_outputs(4470));
    layer1_outputs(4542) <= not(layer0_outputs(895));
    layer1_outputs(4543) <= layer0_outputs(8581);
    layer1_outputs(4544) <= not(layer0_outputs(2235));
    layer1_outputs(4545) <= (layer0_outputs(2364)) and not (layer0_outputs(8777));
    layer1_outputs(4546) <= not(layer0_outputs(10001)) or (layer0_outputs(7006));
    layer1_outputs(4547) <= (layer0_outputs(2825)) and (layer0_outputs(3191));
    layer1_outputs(4548) <= not(layer0_outputs(4410)) or (layer0_outputs(6569));
    layer1_outputs(4549) <= not(layer0_outputs(3911));
    layer1_outputs(4550) <= layer0_outputs(6049);
    layer1_outputs(4551) <= (layer0_outputs(9700)) and not (layer0_outputs(8411));
    layer1_outputs(4552) <= layer0_outputs(9801);
    layer1_outputs(4553) <= not(layer0_outputs(3972));
    layer1_outputs(4554) <= (layer0_outputs(8102)) and (layer0_outputs(5684));
    layer1_outputs(4555) <= layer0_outputs(7868);
    layer1_outputs(4556) <= not(layer0_outputs(4749));
    layer1_outputs(4557) <= not(layer0_outputs(5609));
    layer1_outputs(4558) <= '1';
    layer1_outputs(4559) <= (layer0_outputs(4220)) xor (layer0_outputs(1115));
    layer1_outputs(4560) <= layer0_outputs(430);
    layer1_outputs(4561) <= layer0_outputs(3886);
    layer1_outputs(4562) <= not(layer0_outputs(4722)) or (layer0_outputs(1694));
    layer1_outputs(4563) <= (layer0_outputs(7995)) xor (layer0_outputs(5330));
    layer1_outputs(4564) <= (layer0_outputs(2390)) and not (layer0_outputs(4214));
    layer1_outputs(4565) <= (layer0_outputs(3692)) and not (layer0_outputs(4891));
    layer1_outputs(4566) <= layer0_outputs(9164);
    layer1_outputs(4567) <= (layer0_outputs(5871)) or (layer0_outputs(263));
    layer1_outputs(4568) <= not(layer0_outputs(6685));
    layer1_outputs(4569) <= layer0_outputs(9024);
    layer1_outputs(4570) <= not(layer0_outputs(1442));
    layer1_outputs(4571) <= not(layer0_outputs(1405));
    layer1_outputs(4572) <= layer0_outputs(7478);
    layer1_outputs(4573) <= not((layer0_outputs(10111)) and (layer0_outputs(1582)));
    layer1_outputs(4574) <= not(layer0_outputs(7597));
    layer1_outputs(4575) <= not(layer0_outputs(9168));
    layer1_outputs(4576) <= layer0_outputs(3577);
    layer1_outputs(4577) <= (layer0_outputs(1404)) and not (layer0_outputs(6784));
    layer1_outputs(4578) <= layer0_outputs(4095);
    layer1_outputs(4579) <= not((layer0_outputs(7955)) or (layer0_outputs(4199)));
    layer1_outputs(4580) <= not((layer0_outputs(5709)) and (layer0_outputs(385)));
    layer1_outputs(4581) <= layer0_outputs(9043);
    layer1_outputs(4582) <= layer0_outputs(8358);
    layer1_outputs(4583) <= not((layer0_outputs(1508)) or (layer0_outputs(8378)));
    layer1_outputs(4584) <= layer0_outputs(351);
    layer1_outputs(4585) <= not(layer0_outputs(222));
    layer1_outputs(4586) <= '0';
    layer1_outputs(4587) <= '0';
    layer1_outputs(4588) <= not((layer0_outputs(630)) or (layer0_outputs(2654)));
    layer1_outputs(4589) <= not(layer0_outputs(4548));
    layer1_outputs(4590) <= not((layer0_outputs(9606)) xor (layer0_outputs(7771)));
    layer1_outputs(4591) <= (layer0_outputs(2424)) or (layer0_outputs(9317));
    layer1_outputs(4592) <= not(layer0_outputs(2969));
    layer1_outputs(4593) <= not((layer0_outputs(7120)) or (layer0_outputs(9320)));
    layer1_outputs(4594) <= not(layer0_outputs(5646));
    layer1_outputs(4595) <= not(layer0_outputs(4679));
    layer1_outputs(4596) <= not(layer0_outputs(6329));
    layer1_outputs(4597) <= (layer0_outputs(6508)) and (layer0_outputs(7550));
    layer1_outputs(4598) <= layer0_outputs(628);
    layer1_outputs(4599) <= not((layer0_outputs(1743)) and (layer0_outputs(1951)));
    layer1_outputs(4600) <= not((layer0_outputs(2059)) and (layer0_outputs(6981)));
    layer1_outputs(4601) <= not(layer0_outputs(1939)) or (layer0_outputs(9326));
    layer1_outputs(4602) <= (layer0_outputs(1701)) and not (layer0_outputs(3033));
    layer1_outputs(4603) <= not(layer0_outputs(1810));
    layer1_outputs(4604) <= (layer0_outputs(1463)) and (layer0_outputs(5259));
    layer1_outputs(4605) <= (layer0_outputs(9092)) and (layer0_outputs(8602));
    layer1_outputs(4606) <= not(layer0_outputs(1406));
    layer1_outputs(4607) <= not(layer0_outputs(168)) or (layer0_outputs(5726));
    layer1_outputs(4608) <= layer0_outputs(456);
    layer1_outputs(4609) <= not((layer0_outputs(555)) xor (layer0_outputs(7472)));
    layer1_outputs(4610) <= (layer0_outputs(8026)) and not (layer0_outputs(349));
    layer1_outputs(4611) <= (layer0_outputs(7848)) and not (layer0_outputs(2198));
    layer1_outputs(4612) <= layer0_outputs(6977);
    layer1_outputs(4613) <= (layer0_outputs(3154)) and not (layer0_outputs(3254));
    layer1_outputs(4614) <= layer0_outputs(1352);
    layer1_outputs(4615) <= not(layer0_outputs(5463));
    layer1_outputs(4616) <= not((layer0_outputs(6626)) and (layer0_outputs(5821)));
    layer1_outputs(4617) <= '0';
    layer1_outputs(4618) <= (layer0_outputs(5747)) xor (layer0_outputs(7691));
    layer1_outputs(4619) <= not((layer0_outputs(4150)) xor (layer0_outputs(713)));
    layer1_outputs(4620) <= not((layer0_outputs(8546)) or (layer0_outputs(5752)));
    layer1_outputs(4621) <= not((layer0_outputs(5343)) and (layer0_outputs(7722)));
    layer1_outputs(4622) <= layer0_outputs(2755);
    layer1_outputs(4623) <= not((layer0_outputs(1604)) and (layer0_outputs(1286)));
    layer1_outputs(4624) <= not((layer0_outputs(5414)) and (layer0_outputs(4743)));
    layer1_outputs(4625) <= layer0_outputs(6386);
    layer1_outputs(4626) <= not(layer0_outputs(2181)) or (layer0_outputs(1296));
    layer1_outputs(4627) <= not((layer0_outputs(143)) and (layer0_outputs(5545)));
    layer1_outputs(4628) <= (layer0_outputs(4334)) and not (layer0_outputs(4486));
    layer1_outputs(4629) <= not((layer0_outputs(204)) or (layer0_outputs(7341)));
    layer1_outputs(4630) <= not((layer0_outputs(4472)) or (layer0_outputs(1980)));
    layer1_outputs(4631) <= not((layer0_outputs(3205)) and (layer0_outputs(1155)));
    layer1_outputs(4632) <= (layer0_outputs(2058)) or (layer0_outputs(5162));
    layer1_outputs(4633) <= not(layer0_outputs(514)) or (layer0_outputs(9054));
    layer1_outputs(4634) <= not(layer0_outputs(6763));
    layer1_outputs(4635) <= layer0_outputs(139);
    layer1_outputs(4636) <= (layer0_outputs(428)) xor (layer0_outputs(4599));
    layer1_outputs(4637) <= layer0_outputs(6424);
    layer1_outputs(4638) <= not(layer0_outputs(3247)) or (layer0_outputs(8491));
    layer1_outputs(4639) <= (layer0_outputs(3640)) or (layer0_outputs(8311));
    layer1_outputs(4640) <= not((layer0_outputs(5340)) or (layer0_outputs(2090)));
    layer1_outputs(4641) <= layer0_outputs(4227);
    layer1_outputs(4642) <= (layer0_outputs(962)) xor (layer0_outputs(618));
    layer1_outputs(4643) <= (layer0_outputs(9448)) or (layer0_outputs(3706));
    layer1_outputs(4644) <= not(layer0_outputs(5492)) or (layer0_outputs(5850));
    layer1_outputs(4645) <= not(layer0_outputs(2543)) or (layer0_outputs(3486));
    layer1_outputs(4646) <= (layer0_outputs(7776)) and not (layer0_outputs(7449));
    layer1_outputs(4647) <= '1';
    layer1_outputs(4648) <= not((layer0_outputs(7462)) or (layer0_outputs(620)));
    layer1_outputs(4649) <= (layer0_outputs(9959)) and (layer0_outputs(2271));
    layer1_outputs(4650) <= (layer0_outputs(4975)) and (layer0_outputs(5374));
    layer1_outputs(4651) <= layer0_outputs(7592);
    layer1_outputs(4652) <= not(layer0_outputs(1289));
    layer1_outputs(4653) <= (layer0_outputs(9162)) and not (layer0_outputs(9950));
    layer1_outputs(4654) <= (layer0_outputs(194)) and not (layer0_outputs(4982));
    layer1_outputs(4655) <= (layer0_outputs(1180)) and not (layer0_outputs(7682));
    layer1_outputs(4656) <= layer0_outputs(7951);
    layer1_outputs(4657) <= not((layer0_outputs(4405)) and (layer0_outputs(2467)));
    layer1_outputs(4658) <= not((layer0_outputs(5660)) or (layer0_outputs(1965)));
    layer1_outputs(4659) <= not((layer0_outputs(4996)) xor (layer0_outputs(2864)));
    layer1_outputs(4660) <= (layer0_outputs(131)) and (layer0_outputs(8185));
    layer1_outputs(4661) <= layer0_outputs(4626);
    layer1_outputs(4662) <= not((layer0_outputs(10228)) xor (layer0_outputs(9339)));
    layer1_outputs(4663) <= not(layer0_outputs(4092)) or (layer0_outputs(7391));
    layer1_outputs(4664) <= layer0_outputs(645);
    layer1_outputs(4665) <= (layer0_outputs(9966)) and (layer0_outputs(5808));
    layer1_outputs(4666) <= layer0_outputs(8224);
    layer1_outputs(4667) <= layer0_outputs(6362);
    layer1_outputs(4668) <= not(layer0_outputs(2774)) or (layer0_outputs(3335));
    layer1_outputs(4669) <= not(layer0_outputs(9086)) or (layer0_outputs(4879));
    layer1_outputs(4670) <= layer0_outputs(6320);
    layer1_outputs(4671) <= not((layer0_outputs(3807)) or (layer0_outputs(4338)));
    layer1_outputs(4672) <= layer0_outputs(660);
    layer1_outputs(4673) <= not((layer0_outputs(4706)) xor (layer0_outputs(8459)));
    layer1_outputs(4674) <= not(layer0_outputs(7247));
    layer1_outputs(4675) <= '0';
    layer1_outputs(4676) <= not((layer0_outputs(7386)) or (layer0_outputs(1177)));
    layer1_outputs(4677) <= not(layer0_outputs(4339)) or (layer0_outputs(5689));
    layer1_outputs(4678) <= not(layer0_outputs(5419)) or (layer0_outputs(3053));
    layer1_outputs(4679) <= not(layer0_outputs(849)) or (layer0_outputs(4791));
    layer1_outputs(4680) <= layer0_outputs(1553);
    layer1_outputs(4681) <= layer0_outputs(33);
    layer1_outputs(4682) <= not(layer0_outputs(5762));
    layer1_outputs(4683) <= not(layer0_outputs(1489));
    layer1_outputs(4684) <= (layer0_outputs(2647)) and not (layer0_outputs(4795));
    layer1_outputs(4685) <= not(layer0_outputs(3141));
    layer1_outputs(4686) <= not(layer0_outputs(3422));
    layer1_outputs(4687) <= layer0_outputs(4558);
    layer1_outputs(4688) <= (layer0_outputs(8139)) and not (layer0_outputs(2083));
    layer1_outputs(4689) <= not(layer0_outputs(2715)) or (layer0_outputs(394));
    layer1_outputs(4690) <= not(layer0_outputs(7539));
    layer1_outputs(4691) <= not(layer0_outputs(2291));
    layer1_outputs(4692) <= not((layer0_outputs(7034)) and (layer0_outputs(5976)));
    layer1_outputs(4693) <= not(layer0_outputs(6557));
    layer1_outputs(4694) <= (layer0_outputs(2237)) or (layer0_outputs(2499));
    layer1_outputs(4695) <= (layer0_outputs(3810)) xor (layer0_outputs(6342));
    layer1_outputs(4696) <= (layer0_outputs(4206)) and not (layer0_outputs(7698));
    layer1_outputs(4697) <= not(layer0_outputs(4139)) or (layer0_outputs(2998));
    layer1_outputs(4698) <= not(layer0_outputs(8894)) or (layer0_outputs(8523));
    layer1_outputs(4699) <= not(layer0_outputs(5577));
    layer1_outputs(4700) <= layer0_outputs(9664);
    layer1_outputs(4701) <= not((layer0_outputs(5686)) xor (layer0_outputs(10018)));
    layer1_outputs(4702) <= not(layer0_outputs(9479)) or (layer0_outputs(430));
    layer1_outputs(4703) <= (layer0_outputs(2365)) and (layer0_outputs(1167));
    layer1_outputs(4704) <= (layer0_outputs(6918)) and not (layer0_outputs(7028));
    layer1_outputs(4705) <= not((layer0_outputs(7603)) xor (layer0_outputs(9191)));
    layer1_outputs(4706) <= (layer0_outputs(5357)) or (layer0_outputs(4829));
    layer1_outputs(4707) <= not(layer0_outputs(3105)) or (layer0_outputs(4809));
    layer1_outputs(4708) <= layer0_outputs(624);
    layer1_outputs(4709) <= not(layer0_outputs(295));
    layer1_outputs(4710) <= not(layer0_outputs(2831));
    layer1_outputs(4711) <= not(layer0_outputs(6516));
    layer1_outputs(4712) <= layer0_outputs(4308);
    layer1_outputs(4713) <= (layer0_outputs(6658)) and (layer0_outputs(749));
    layer1_outputs(4714) <= not((layer0_outputs(4006)) and (layer0_outputs(1632)));
    layer1_outputs(4715) <= layer0_outputs(2490);
    layer1_outputs(4716) <= layer0_outputs(8107);
    layer1_outputs(4717) <= not(layer0_outputs(2008));
    layer1_outputs(4718) <= not(layer0_outputs(9370)) or (layer0_outputs(438));
    layer1_outputs(4719) <= (layer0_outputs(6148)) xor (layer0_outputs(9655));
    layer1_outputs(4720) <= not(layer0_outputs(1169)) or (layer0_outputs(6138));
    layer1_outputs(4721) <= not(layer0_outputs(2475));
    layer1_outputs(4722) <= not(layer0_outputs(4944));
    layer1_outputs(4723) <= not(layer0_outputs(5892)) or (layer0_outputs(237));
    layer1_outputs(4724) <= (layer0_outputs(1600)) and (layer0_outputs(7030));
    layer1_outputs(4725) <= layer0_outputs(5391);
    layer1_outputs(4726) <= (layer0_outputs(4500)) or (layer0_outputs(5061));
    layer1_outputs(4727) <= not(layer0_outputs(5115));
    layer1_outputs(4728) <= (layer0_outputs(471)) or (layer0_outputs(9044));
    layer1_outputs(4729) <= (layer0_outputs(7776)) or (layer0_outputs(5915));
    layer1_outputs(4730) <= not(layer0_outputs(509));
    layer1_outputs(4731) <= (layer0_outputs(1066)) or (layer0_outputs(8327));
    layer1_outputs(4732) <= not((layer0_outputs(6638)) xor (layer0_outputs(4558)));
    layer1_outputs(4733) <= layer0_outputs(9278);
    layer1_outputs(4734) <= not(layer0_outputs(6713)) or (layer0_outputs(5979));
    layer1_outputs(4735) <= not(layer0_outputs(926));
    layer1_outputs(4736) <= (layer0_outputs(2128)) and not (layer0_outputs(8016));
    layer1_outputs(4737) <= layer0_outputs(9282);
    layer1_outputs(4738) <= layer0_outputs(7922);
    layer1_outputs(4739) <= layer0_outputs(6519);
    layer1_outputs(4740) <= (layer0_outputs(6984)) xor (layer0_outputs(7277));
    layer1_outputs(4741) <= not((layer0_outputs(9197)) or (layer0_outputs(6039)));
    layer1_outputs(4742) <= not(layer0_outputs(34));
    layer1_outputs(4743) <= not(layer0_outputs(2196));
    layer1_outputs(4744) <= not((layer0_outputs(7875)) xor (layer0_outputs(2961)));
    layer1_outputs(4745) <= layer0_outputs(9618);
    layer1_outputs(4746) <= not(layer0_outputs(5904)) or (layer0_outputs(976));
    layer1_outputs(4747) <= (layer0_outputs(9398)) and (layer0_outputs(6484));
    layer1_outputs(4748) <= (layer0_outputs(5305)) and not (layer0_outputs(628));
    layer1_outputs(4749) <= not((layer0_outputs(5877)) or (layer0_outputs(5186)));
    layer1_outputs(4750) <= not(layer0_outputs(6169));
    layer1_outputs(4751) <= not((layer0_outputs(9385)) or (layer0_outputs(9856)));
    layer1_outputs(4752) <= not(layer0_outputs(5272));
    layer1_outputs(4753) <= layer0_outputs(9797);
    layer1_outputs(4754) <= (layer0_outputs(5203)) and not (layer0_outputs(5350));
    layer1_outputs(4755) <= not(layer0_outputs(9786)) or (layer0_outputs(2433));
    layer1_outputs(4756) <= not((layer0_outputs(6344)) xor (layer0_outputs(662)));
    layer1_outputs(4757) <= (layer0_outputs(6943)) xor (layer0_outputs(10027));
    layer1_outputs(4758) <= layer0_outputs(7518);
    layer1_outputs(4759) <= layer0_outputs(3687);
    layer1_outputs(4760) <= not((layer0_outputs(8574)) or (layer0_outputs(1465)));
    layer1_outputs(4761) <= (layer0_outputs(6735)) and (layer0_outputs(3825));
    layer1_outputs(4762) <= not(layer0_outputs(1180)) or (layer0_outputs(8856));
    layer1_outputs(4763) <= (layer0_outputs(2709)) and not (layer0_outputs(1736));
    layer1_outputs(4764) <= not(layer0_outputs(3780));
    layer1_outputs(4765) <= not((layer0_outputs(6491)) and (layer0_outputs(2178)));
    layer1_outputs(4766) <= not(layer0_outputs(2070)) or (layer0_outputs(8733));
    layer1_outputs(4767) <= layer0_outputs(8927);
    layer1_outputs(4768) <= not(layer0_outputs(9390)) or (layer0_outputs(9480));
    layer1_outputs(4769) <= not(layer0_outputs(4304));
    layer1_outputs(4770) <= (layer0_outputs(9458)) and not (layer0_outputs(703));
    layer1_outputs(4771) <= layer0_outputs(8630);
    layer1_outputs(4772) <= not(layer0_outputs(3769));
    layer1_outputs(4773) <= layer0_outputs(1628);
    layer1_outputs(4774) <= not((layer0_outputs(112)) or (layer0_outputs(3594)));
    layer1_outputs(4775) <= (layer0_outputs(1641)) and not (layer0_outputs(5195));
    layer1_outputs(4776) <= not((layer0_outputs(1940)) or (layer0_outputs(6762)));
    layer1_outputs(4777) <= not(layer0_outputs(2797));
    layer1_outputs(4778) <= not(layer0_outputs(245));
    layer1_outputs(4779) <= (layer0_outputs(9473)) and not (layer0_outputs(3353));
    layer1_outputs(4780) <= layer0_outputs(5594);
    layer1_outputs(4781) <= not(layer0_outputs(9333));
    layer1_outputs(4782) <= not(layer0_outputs(7636));
    layer1_outputs(4783) <= (layer0_outputs(973)) and not (layer0_outputs(3562));
    layer1_outputs(4784) <= not((layer0_outputs(10116)) xor (layer0_outputs(5277)));
    layer1_outputs(4785) <= not((layer0_outputs(1361)) and (layer0_outputs(10177)));
    layer1_outputs(4786) <= layer0_outputs(910);
    layer1_outputs(4787) <= '0';
    layer1_outputs(4788) <= not((layer0_outputs(4340)) or (layer0_outputs(4248)));
    layer1_outputs(4789) <= '1';
    layer1_outputs(4790) <= layer0_outputs(4552);
    layer1_outputs(4791) <= (layer0_outputs(3565)) xor (layer0_outputs(6539));
    layer1_outputs(4792) <= (layer0_outputs(6049)) xor (layer0_outputs(5292));
    layer1_outputs(4793) <= layer0_outputs(5502);
    layer1_outputs(4794) <= (layer0_outputs(10096)) and (layer0_outputs(10229));
    layer1_outputs(4795) <= not(layer0_outputs(5315)) or (layer0_outputs(9956));
    layer1_outputs(4796) <= '1';
    layer1_outputs(4797) <= layer0_outputs(3309);
    layer1_outputs(4798) <= (layer0_outputs(7785)) xor (layer0_outputs(8072));
    layer1_outputs(4799) <= (layer0_outputs(8513)) and not (layer0_outputs(4423));
    layer1_outputs(4800) <= '1';
    layer1_outputs(4801) <= layer0_outputs(6189);
    layer1_outputs(4802) <= not(layer0_outputs(1715));
    layer1_outputs(4803) <= (layer0_outputs(2379)) and not (layer0_outputs(5839));
    layer1_outputs(4804) <= layer0_outputs(8715);
    layer1_outputs(4805) <= not(layer0_outputs(9193));
    layer1_outputs(4806) <= not((layer0_outputs(7655)) xor (layer0_outputs(7772)));
    layer1_outputs(4807) <= '0';
    layer1_outputs(4808) <= not((layer0_outputs(5900)) and (layer0_outputs(1318)));
    layer1_outputs(4809) <= (layer0_outputs(1163)) and not (layer0_outputs(6295));
    layer1_outputs(4810) <= not(layer0_outputs(4716));
    layer1_outputs(4811) <= not(layer0_outputs(3654)) or (layer0_outputs(5561));
    layer1_outputs(4812) <= layer0_outputs(8225);
    layer1_outputs(4813) <= (layer0_outputs(7106)) and not (layer0_outputs(643));
    layer1_outputs(4814) <= (layer0_outputs(7311)) or (layer0_outputs(2152));
    layer1_outputs(4815) <= not(layer0_outputs(7673));
    layer1_outputs(4816) <= (layer0_outputs(4969)) or (layer0_outputs(7302));
    layer1_outputs(4817) <= not((layer0_outputs(5064)) and (layer0_outputs(564)));
    layer1_outputs(4818) <= not(layer0_outputs(867)) or (layer0_outputs(2800));
    layer1_outputs(4819) <= layer0_outputs(5194);
    layer1_outputs(4820) <= (layer0_outputs(905)) or (layer0_outputs(7265));
    layer1_outputs(4821) <= not(layer0_outputs(7243)) or (layer0_outputs(5152));
    layer1_outputs(4822) <= not((layer0_outputs(3988)) or (layer0_outputs(2080)));
    layer1_outputs(4823) <= '0';
    layer1_outputs(4824) <= (layer0_outputs(4048)) or (layer0_outputs(9428));
    layer1_outputs(4825) <= not(layer0_outputs(6634));
    layer1_outputs(4826) <= (layer0_outputs(7574)) or (layer0_outputs(2776));
    layer1_outputs(4827) <= layer0_outputs(6688);
    layer1_outputs(4828) <= not(layer0_outputs(4132));
    layer1_outputs(4829) <= not(layer0_outputs(5431));
    layer1_outputs(4830) <= not(layer0_outputs(8308)) or (layer0_outputs(3242));
    layer1_outputs(4831) <= not(layer0_outputs(6425)) or (layer0_outputs(7684));
    layer1_outputs(4832) <= (layer0_outputs(2129)) and not (layer0_outputs(9890));
    layer1_outputs(4833) <= layer0_outputs(4837);
    layer1_outputs(4834) <= layer0_outputs(6630);
    layer1_outputs(4835) <= not((layer0_outputs(4788)) and (layer0_outputs(6194)));
    layer1_outputs(4836) <= not(layer0_outputs(3764)) or (layer0_outputs(2527));
    layer1_outputs(4837) <= not(layer0_outputs(1843));
    layer1_outputs(4838) <= not(layer0_outputs(309)) or (layer0_outputs(8783));
    layer1_outputs(4839) <= not(layer0_outputs(6631));
    layer1_outputs(4840) <= not(layer0_outputs(7008));
    layer1_outputs(4841) <= not(layer0_outputs(1301)) or (layer0_outputs(3243));
    layer1_outputs(4842) <= not((layer0_outputs(6903)) or (layer0_outputs(9237)));
    layer1_outputs(4843) <= '0';
    layer1_outputs(4844) <= not(layer0_outputs(3524));
    layer1_outputs(4845) <= layer0_outputs(4178);
    layer1_outputs(4846) <= not((layer0_outputs(7808)) or (layer0_outputs(2837)));
    layer1_outputs(4847) <= layer0_outputs(7209);
    layer1_outputs(4848) <= not(layer0_outputs(6043));
    layer1_outputs(4849) <= not(layer0_outputs(857));
    layer1_outputs(4850) <= (layer0_outputs(2021)) or (layer0_outputs(211));
    layer1_outputs(4851) <= not(layer0_outputs(28));
    layer1_outputs(4852) <= (layer0_outputs(6704)) and (layer0_outputs(5571));
    layer1_outputs(4853) <= layer0_outputs(9833);
    layer1_outputs(4854) <= not(layer0_outputs(2611));
    layer1_outputs(4855) <= (layer0_outputs(2127)) and not (layer0_outputs(2345));
    layer1_outputs(4856) <= not((layer0_outputs(6221)) or (layer0_outputs(6726)));
    layer1_outputs(4857) <= not((layer0_outputs(5021)) and (layer0_outputs(958)));
    layer1_outputs(4858) <= not(layer0_outputs(2947)) or (layer0_outputs(6018));
    layer1_outputs(4859) <= not((layer0_outputs(9556)) xor (layer0_outputs(10198)));
    layer1_outputs(4860) <= (layer0_outputs(3999)) and not (layer0_outputs(10178));
    layer1_outputs(4861) <= (layer0_outputs(8498)) xor (layer0_outputs(4177));
    layer1_outputs(4862) <= not((layer0_outputs(7599)) and (layer0_outputs(9833)));
    layer1_outputs(4863) <= layer0_outputs(6577);
    layer1_outputs(4864) <= not(layer0_outputs(8090)) or (layer0_outputs(8148));
    layer1_outputs(4865) <= (layer0_outputs(6118)) and (layer0_outputs(8304));
    layer1_outputs(4866) <= layer0_outputs(8877);
    layer1_outputs(4867) <= (layer0_outputs(167)) and not (layer0_outputs(4193));
    layer1_outputs(4868) <= not(layer0_outputs(7760)) or (layer0_outputs(9394));
    layer1_outputs(4869) <= '0';
    layer1_outputs(4870) <= (layer0_outputs(8191)) and not (layer0_outputs(8467));
    layer1_outputs(4871) <= layer0_outputs(7446);
    layer1_outputs(4872) <= not(layer0_outputs(5411));
    layer1_outputs(4873) <= '1';
    layer1_outputs(4874) <= layer0_outputs(2090);
    layer1_outputs(4875) <= not(layer0_outputs(3094)) or (layer0_outputs(9099));
    layer1_outputs(4876) <= (layer0_outputs(7001)) and not (layer0_outputs(2277));
    layer1_outputs(4877) <= layer0_outputs(9159);
    layer1_outputs(4878) <= (layer0_outputs(4330)) and not (layer0_outputs(9242));
    layer1_outputs(4879) <= (layer0_outputs(7363)) xor (layer0_outputs(4565));
    layer1_outputs(4880) <= (layer0_outputs(8247)) xor (layer0_outputs(9741));
    layer1_outputs(4881) <= (layer0_outputs(49)) and not (layer0_outputs(7978));
    layer1_outputs(4882) <= not(layer0_outputs(3185)) or (layer0_outputs(5556));
    layer1_outputs(4883) <= (layer0_outputs(724)) xor (layer0_outputs(4972));
    layer1_outputs(4884) <= layer0_outputs(2329);
    layer1_outputs(4885) <= (layer0_outputs(9828)) and not (layer0_outputs(9785));
    layer1_outputs(4886) <= not(layer0_outputs(8984)) or (layer0_outputs(5024));
    layer1_outputs(4887) <= not((layer0_outputs(6738)) and (layer0_outputs(4231)));
    layer1_outputs(4888) <= (layer0_outputs(107)) and not (layer0_outputs(4892));
    layer1_outputs(4889) <= layer0_outputs(6623);
    layer1_outputs(4890) <= (layer0_outputs(9740)) xor (layer0_outputs(1663));
    layer1_outputs(4891) <= not(layer0_outputs(5797));
    layer1_outputs(4892) <= (layer0_outputs(2944)) xor (layer0_outputs(2944));
    layer1_outputs(4893) <= not((layer0_outputs(7844)) or (layer0_outputs(2846)));
    layer1_outputs(4894) <= (layer0_outputs(8155)) or (layer0_outputs(2132));
    layer1_outputs(4895) <= not(layer0_outputs(10069));
    layer1_outputs(4896) <= not((layer0_outputs(4379)) xor (layer0_outputs(1548)));
    layer1_outputs(4897) <= not((layer0_outputs(4715)) and (layer0_outputs(8597)));
    layer1_outputs(4898) <= not(layer0_outputs(4014));
    layer1_outputs(4899) <= not((layer0_outputs(1436)) and (layer0_outputs(1242)));
    layer1_outputs(4900) <= layer0_outputs(8783);
    layer1_outputs(4901) <= not(layer0_outputs(3157)) or (layer0_outputs(7394));
    layer1_outputs(4902) <= layer0_outputs(5554);
    layer1_outputs(4903) <= (layer0_outputs(7990)) and not (layer0_outputs(5969));
    layer1_outputs(4904) <= not((layer0_outputs(9944)) xor (layer0_outputs(5926)));
    layer1_outputs(4905) <= not(layer0_outputs(4968));
    layer1_outputs(4906) <= not((layer0_outputs(946)) or (layer0_outputs(6394)));
    layer1_outputs(4907) <= (layer0_outputs(1582)) and not (layer0_outputs(1023));
    layer1_outputs(4908) <= not((layer0_outputs(10040)) xor (layer0_outputs(1119)));
    layer1_outputs(4909) <= (layer0_outputs(909)) and not (layer0_outputs(8031));
    layer1_outputs(4910) <= not(layer0_outputs(8655)) or (layer0_outputs(2250));
    layer1_outputs(4911) <= layer0_outputs(2681);
    layer1_outputs(4912) <= (layer0_outputs(7260)) and not (layer0_outputs(64));
    layer1_outputs(4913) <= not((layer0_outputs(3957)) and (layer0_outputs(3117)));
    layer1_outputs(4914) <= not(layer0_outputs(8056));
    layer1_outputs(4915) <= not(layer0_outputs(9128));
    layer1_outputs(4916) <= (layer0_outputs(3035)) and (layer0_outputs(5316));
    layer1_outputs(4917) <= not(layer0_outputs(4472)) or (layer0_outputs(9401));
    layer1_outputs(4918) <= layer0_outputs(1186);
    layer1_outputs(4919) <= not((layer0_outputs(3274)) and (layer0_outputs(4985)));
    layer1_outputs(4920) <= (layer0_outputs(328)) and not (layer0_outputs(6790));
    layer1_outputs(4921) <= (layer0_outputs(3520)) and not (layer0_outputs(7113));
    layer1_outputs(4922) <= not(layer0_outputs(203));
    layer1_outputs(4923) <= not((layer0_outputs(3573)) xor (layer0_outputs(2429)));
    layer1_outputs(4924) <= '1';
    layer1_outputs(4925) <= not(layer0_outputs(1966));
    layer1_outputs(4926) <= not(layer0_outputs(1870));
    layer1_outputs(4927) <= (layer0_outputs(9066)) and (layer0_outputs(5402));
    layer1_outputs(4928) <= not(layer0_outputs(2018));
    layer1_outputs(4929) <= not((layer0_outputs(4973)) xor (layer0_outputs(9596)));
    layer1_outputs(4930) <= (layer0_outputs(9733)) and not (layer0_outputs(7563));
    layer1_outputs(4931) <= (layer0_outputs(8677)) and not (layer0_outputs(9353));
    layer1_outputs(4932) <= layer0_outputs(1261);
    layer1_outputs(4933) <= '0';
    layer1_outputs(4934) <= not((layer0_outputs(1398)) xor (layer0_outputs(6760)));
    layer1_outputs(4935) <= not((layer0_outputs(9298)) or (layer0_outputs(6731)));
    layer1_outputs(4936) <= (layer0_outputs(1003)) and not (layer0_outputs(7482));
    layer1_outputs(4937) <= not((layer0_outputs(3680)) and (layer0_outputs(3927)));
    layer1_outputs(4938) <= not((layer0_outputs(1872)) and (layer0_outputs(6274)));
    layer1_outputs(4939) <= not((layer0_outputs(3142)) or (layer0_outputs(9646)));
    layer1_outputs(4940) <= not(layer0_outputs(1742));
    layer1_outputs(4941) <= layer0_outputs(3453);
    layer1_outputs(4942) <= not(layer0_outputs(8836));
    layer1_outputs(4943) <= not(layer0_outputs(2299));
    layer1_outputs(4944) <= layer0_outputs(3220);
    layer1_outputs(4945) <= not(layer0_outputs(9685));
    layer1_outputs(4946) <= not(layer0_outputs(8628));
    layer1_outputs(4947) <= layer0_outputs(9196);
    layer1_outputs(4948) <= not(layer0_outputs(6476));
    layer1_outputs(4949) <= (layer0_outputs(4601)) or (layer0_outputs(5693));
    layer1_outputs(4950) <= (layer0_outputs(2075)) and not (layer0_outputs(10029));
    layer1_outputs(4951) <= (layer0_outputs(3472)) and not (layer0_outputs(4284));
    layer1_outputs(4952) <= '0';
    layer1_outputs(4953) <= not(layer0_outputs(7111)) or (layer0_outputs(2686));
    layer1_outputs(4954) <= not((layer0_outputs(9481)) or (layer0_outputs(3799)));
    layer1_outputs(4955) <= (layer0_outputs(4819)) or (layer0_outputs(7548));
    layer1_outputs(4956) <= (layer0_outputs(7327)) and not (layer0_outputs(2353));
    layer1_outputs(4957) <= not((layer0_outputs(3771)) xor (layer0_outputs(1615)));
    layer1_outputs(4958) <= not((layer0_outputs(2706)) xor (layer0_outputs(8410)));
    layer1_outputs(4959) <= (layer0_outputs(5879)) and (layer0_outputs(9593));
    layer1_outputs(4960) <= (layer0_outputs(2219)) or (layer0_outputs(1762));
    layer1_outputs(4961) <= not((layer0_outputs(8937)) and (layer0_outputs(5484)));
    layer1_outputs(4962) <= (layer0_outputs(1905)) and (layer0_outputs(95));
    layer1_outputs(4963) <= (layer0_outputs(1354)) and not (layer0_outputs(5349));
    layer1_outputs(4964) <= not(layer0_outputs(163));
    layer1_outputs(4965) <= not(layer0_outputs(1856));
    layer1_outputs(4966) <= not(layer0_outputs(7422));
    layer1_outputs(4967) <= not(layer0_outputs(1223));
    layer1_outputs(4968) <= (layer0_outputs(2331)) and not (layer0_outputs(725));
    layer1_outputs(4969) <= not(layer0_outputs(3918));
    layer1_outputs(4970) <= not(layer0_outputs(5771));
    layer1_outputs(4971) <= layer0_outputs(7953);
    layer1_outputs(4972) <= not(layer0_outputs(2000));
    layer1_outputs(4973) <= layer0_outputs(5058);
    layer1_outputs(4974) <= not(layer0_outputs(6901));
    layer1_outputs(4975) <= layer0_outputs(10104);
    layer1_outputs(4976) <= (layer0_outputs(2876)) or (layer0_outputs(5358));
    layer1_outputs(4977) <= (layer0_outputs(10107)) or (layer0_outputs(8048));
    layer1_outputs(4978) <= layer0_outputs(6230);
    layer1_outputs(4979) <= not((layer0_outputs(1731)) and (layer0_outputs(6972)));
    layer1_outputs(4980) <= not(layer0_outputs(6651));
    layer1_outputs(4981) <= not(layer0_outputs(3997));
    layer1_outputs(4982) <= layer0_outputs(3023);
    layer1_outputs(4983) <= not(layer0_outputs(5286)) or (layer0_outputs(2259));
    layer1_outputs(4984) <= not(layer0_outputs(9733));
    layer1_outputs(4985) <= (layer0_outputs(3798)) and not (layer0_outputs(7333));
    layer1_outputs(4986) <= (layer0_outputs(3887)) and not (layer0_outputs(8089));
    layer1_outputs(4987) <= not((layer0_outputs(106)) or (layer0_outputs(8929)));
    layer1_outputs(4988) <= not(layer0_outputs(8510));
    layer1_outputs(4989) <= not(layer0_outputs(10034)) or (layer0_outputs(7564));
    layer1_outputs(4990) <= not((layer0_outputs(8148)) xor (layer0_outputs(6579)));
    layer1_outputs(4991) <= (layer0_outputs(3377)) or (layer0_outputs(2450));
    layer1_outputs(4992) <= layer0_outputs(8077);
    layer1_outputs(4993) <= not(layer0_outputs(6538));
    layer1_outputs(4994) <= not((layer0_outputs(2287)) xor (layer0_outputs(8043)));
    layer1_outputs(4995) <= not(layer0_outputs(7384)) or (layer0_outputs(1228));
    layer1_outputs(4996) <= not(layer0_outputs(1264)) or (layer0_outputs(4659));
    layer1_outputs(4997) <= not(layer0_outputs(2957)) or (layer0_outputs(987));
    layer1_outputs(4998) <= layer0_outputs(5541);
    layer1_outputs(4999) <= (layer0_outputs(6850)) or (layer0_outputs(6696));
    layer1_outputs(5000) <= (layer0_outputs(4329)) xor (layer0_outputs(3664));
    layer1_outputs(5001) <= not(layer0_outputs(1052));
    layer1_outputs(5002) <= not(layer0_outputs(4865)) or (layer0_outputs(526));
    layer1_outputs(5003) <= not(layer0_outputs(9883));
    layer1_outputs(5004) <= (layer0_outputs(8900)) and not (layer0_outputs(3872));
    layer1_outputs(5005) <= layer0_outputs(1719);
    layer1_outputs(5006) <= not(layer0_outputs(7777)) or (layer0_outputs(3272));
    layer1_outputs(5007) <= (layer0_outputs(4818)) xor (layer0_outputs(2687));
    layer1_outputs(5008) <= not(layer0_outputs(8532));
    layer1_outputs(5009) <= not((layer0_outputs(3178)) xor (layer0_outputs(6528)));
    layer1_outputs(5010) <= (layer0_outputs(7559)) and not (layer0_outputs(147));
    layer1_outputs(5011) <= not((layer0_outputs(7879)) and (layer0_outputs(2796)));
    layer1_outputs(5012) <= not(layer0_outputs(9838)) or (layer0_outputs(3854));
    layer1_outputs(5013) <= (layer0_outputs(4600)) and not (layer0_outputs(6495));
    layer1_outputs(5014) <= '1';
    layer1_outputs(5015) <= layer0_outputs(6353);
    layer1_outputs(5016) <= not((layer0_outputs(2861)) or (layer0_outputs(566)));
    layer1_outputs(5017) <= not(layer0_outputs(5996));
    layer1_outputs(5018) <= not(layer0_outputs(8773));
    layer1_outputs(5019) <= (layer0_outputs(8982)) and (layer0_outputs(3738));
    layer1_outputs(5020) <= layer0_outputs(5226);
    layer1_outputs(5021) <= (layer0_outputs(9935)) or (layer0_outputs(6124));
    layer1_outputs(5022) <= (layer0_outputs(7883)) and not (layer0_outputs(7133));
    layer1_outputs(5023) <= (layer0_outputs(2171)) or (layer0_outputs(8375));
    layer1_outputs(5024) <= not(layer0_outputs(511));
    layer1_outputs(5025) <= not((layer0_outputs(4219)) xor (layer0_outputs(8542)));
    layer1_outputs(5026) <= (layer0_outputs(3340)) and not (layer0_outputs(2691));
    layer1_outputs(5027) <= not(layer0_outputs(2057)) or (layer0_outputs(5695));
    layer1_outputs(5028) <= (layer0_outputs(1372)) or (layer0_outputs(108));
    layer1_outputs(5029) <= layer0_outputs(7429);
    layer1_outputs(5030) <= not((layer0_outputs(10051)) or (layer0_outputs(5343)));
    layer1_outputs(5031) <= layer0_outputs(6560);
    layer1_outputs(5032) <= (layer0_outputs(9045)) xor (layer0_outputs(7192));
    layer1_outputs(5033) <= not(layer0_outputs(5677));
    layer1_outputs(5034) <= not((layer0_outputs(4657)) xor (layer0_outputs(1625)));
    layer1_outputs(5035) <= layer0_outputs(5579);
    layer1_outputs(5036) <= layer0_outputs(8447);
    layer1_outputs(5037) <= not((layer0_outputs(5099)) and (layer0_outputs(1105)));
    layer1_outputs(5038) <= not(layer0_outputs(1503));
    layer1_outputs(5039) <= not(layer0_outputs(1870));
    layer1_outputs(5040) <= not(layer0_outputs(6897));
    layer1_outputs(5041) <= not((layer0_outputs(9370)) xor (layer0_outputs(9699)));
    layer1_outputs(5042) <= (layer0_outputs(4434)) and not (layer0_outputs(623));
    layer1_outputs(5043) <= not((layer0_outputs(7897)) xor (layer0_outputs(9084)));
    layer1_outputs(5044) <= (layer0_outputs(4907)) and not (layer0_outputs(8478));
    layer1_outputs(5045) <= not((layer0_outputs(8779)) xor (layer0_outputs(4750)));
    layer1_outputs(5046) <= (layer0_outputs(6944)) and not (layer0_outputs(6437));
    layer1_outputs(5047) <= layer0_outputs(4996);
    layer1_outputs(5048) <= not(layer0_outputs(5667)) or (layer0_outputs(9760));
    layer1_outputs(5049) <= (layer0_outputs(5593)) and (layer0_outputs(10001));
    layer1_outputs(5050) <= (layer0_outputs(448)) and not (layer0_outputs(8706));
    layer1_outputs(5051) <= '0';
    layer1_outputs(5052) <= (layer0_outputs(237)) xor (layer0_outputs(4741));
    layer1_outputs(5053) <= layer0_outputs(5532);
    layer1_outputs(5054) <= (layer0_outputs(5987)) and not (layer0_outputs(5352));
    layer1_outputs(5055) <= not(layer0_outputs(8918));
    layer1_outputs(5056) <= (layer0_outputs(9542)) and (layer0_outputs(2032));
    layer1_outputs(5057) <= not((layer0_outputs(4955)) xor (layer0_outputs(4950)));
    layer1_outputs(5058) <= (layer0_outputs(7568)) and not (layer0_outputs(772));
    layer1_outputs(5059) <= layer0_outputs(5375);
    layer1_outputs(5060) <= (layer0_outputs(6735)) and (layer0_outputs(8806));
    layer1_outputs(5061) <= (layer0_outputs(4862)) and (layer0_outputs(3271));
    layer1_outputs(5062) <= layer0_outputs(6639);
    layer1_outputs(5063) <= not(layer0_outputs(9005));
    layer1_outputs(5064) <= (layer0_outputs(7457)) or (layer0_outputs(7608));
    layer1_outputs(5065) <= layer0_outputs(3498);
    layer1_outputs(5066) <= not((layer0_outputs(8804)) xor (layer0_outputs(8854)));
    layer1_outputs(5067) <= not(layer0_outputs(4098));
    layer1_outputs(5068) <= not(layer0_outputs(9963));
    layer1_outputs(5069) <= not((layer0_outputs(8464)) and (layer0_outputs(6248)));
    layer1_outputs(5070) <= not(layer0_outputs(8416));
    layer1_outputs(5071) <= not(layer0_outputs(9553));
    layer1_outputs(5072) <= (layer0_outputs(900)) and (layer0_outputs(2695));
    layer1_outputs(5073) <= layer0_outputs(7338);
    layer1_outputs(5074) <= (layer0_outputs(1407)) and (layer0_outputs(7614));
    layer1_outputs(5075) <= not(layer0_outputs(9449));
    layer1_outputs(5076) <= not(layer0_outputs(5882));
    layer1_outputs(5077) <= layer0_outputs(4825);
    layer1_outputs(5078) <= not(layer0_outputs(1078));
    layer1_outputs(5079) <= (layer0_outputs(7765)) xor (layer0_outputs(8454));
    layer1_outputs(5080) <= (layer0_outputs(3395)) or (layer0_outputs(1807));
    layer1_outputs(5081) <= layer0_outputs(6410);
    layer1_outputs(5082) <= layer0_outputs(1249);
    layer1_outputs(5083) <= not((layer0_outputs(761)) and (layer0_outputs(1835)));
    layer1_outputs(5084) <= not(layer0_outputs(8896)) or (layer0_outputs(10213));
    layer1_outputs(5085) <= not(layer0_outputs(6201)) or (layer0_outputs(6577));
    layer1_outputs(5086) <= not((layer0_outputs(8625)) and (layer0_outputs(10046)));
    layer1_outputs(5087) <= (layer0_outputs(2042)) xor (layer0_outputs(1686));
    layer1_outputs(5088) <= (layer0_outputs(3261)) and not (layer0_outputs(8989));
    layer1_outputs(5089) <= layer0_outputs(1842);
    layer1_outputs(5090) <= (layer0_outputs(6919)) or (layer0_outputs(6176));
    layer1_outputs(5091) <= not((layer0_outputs(223)) or (layer0_outputs(23)));
    layer1_outputs(5092) <= (layer0_outputs(831)) and not (layer0_outputs(6376));
    layer1_outputs(5093) <= layer0_outputs(817);
    layer1_outputs(5094) <= not(layer0_outputs(6040));
    layer1_outputs(5095) <= not(layer0_outputs(2481));
    layer1_outputs(5096) <= (layer0_outputs(5073)) xor (layer0_outputs(1657));
    layer1_outputs(5097) <= (layer0_outputs(8796)) or (layer0_outputs(3070));
    layer1_outputs(5098) <= (layer0_outputs(1166)) or (layer0_outputs(9341));
    layer1_outputs(5099) <= not((layer0_outputs(7970)) and (layer0_outputs(6856)));
    layer1_outputs(5100) <= '0';
    layer1_outputs(5101) <= layer0_outputs(4606);
    layer1_outputs(5102) <= (layer0_outputs(10201)) or (layer0_outputs(8577));
    layer1_outputs(5103) <= not(layer0_outputs(4354));
    layer1_outputs(5104) <= layer0_outputs(1990);
    layer1_outputs(5105) <= (layer0_outputs(7506)) and (layer0_outputs(6506));
    layer1_outputs(5106) <= not((layer0_outputs(4036)) and (layer0_outputs(2476)));
    layer1_outputs(5107) <= not(layer0_outputs(450));
    layer1_outputs(5108) <= not((layer0_outputs(2547)) and (layer0_outputs(8566)));
    layer1_outputs(5109) <= layer0_outputs(261);
    layer1_outputs(5110) <= layer0_outputs(7819);
    layer1_outputs(5111) <= layer0_outputs(3103);
    layer1_outputs(5112) <= not(layer0_outputs(8213));
    layer1_outputs(5113) <= not((layer0_outputs(3988)) and (layer0_outputs(3232)));
    layer1_outputs(5114) <= not((layer0_outputs(1637)) xor (layer0_outputs(3500)));
    layer1_outputs(5115) <= not((layer0_outputs(800)) or (layer0_outputs(7857)));
    layer1_outputs(5116) <= not((layer0_outputs(7026)) or (layer0_outputs(8852)));
    layer1_outputs(5117) <= not((layer0_outputs(1724)) xor (layer0_outputs(2692)));
    layer1_outputs(5118) <= not((layer0_outputs(5680)) or (layer0_outputs(3954)));
    layer1_outputs(5119) <= (layer0_outputs(10050)) and not (layer0_outputs(3371));
    layer1_outputs(5120) <= not(layer0_outputs(2908)) or (layer0_outputs(523));
    layer1_outputs(5121) <= not(layer0_outputs(5476));
    layer1_outputs(5122) <= '1';
    layer1_outputs(5123) <= not(layer0_outputs(6882));
    layer1_outputs(5124) <= layer0_outputs(2713);
    layer1_outputs(5125) <= layer0_outputs(1996);
    layer1_outputs(5126) <= (layer0_outputs(9294)) or (layer0_outputs(5041));
    layer1_outputs(5127) <= not((layer0_outputs(347)) xor (layer0_outputs(2321)));
    layer1_outputs(5128) <= (layer0_outputs(748)) xor (layer0_outputs(9172));
    layer1_outputs(5129) <= layer0_outputs(3543);
    layer1_outputs(5130) <= not(layer0_outputs(4343));
    layer1_outputs(5131) <= not((layer0_outputs(4687)) or (layer0_outputs(4815)));
    layer1_outputs(5132) <= (layer0_outputs(9457)) and (layer0_outputs(2323));
    layer1_outputs(5133) <= (layer0_outputs(3435)) and not (layer0_outputs(2162));
    layer1_outputs(5134) <= (layer0_outputs(3783)) and not (layer0_outputs(741));
    layer1_outputs(5135) <= not(layer0_outputs(2708)) or (layer0_outputs(7870));
    layer1_outputs(5136) <= '0';
    layer1_outputs(5137) <= (layer0_outputs(5602)) and not (layer0_outputs(8714));
    layer1_outputs(5138) <= (layer0_outputs(2100)) and (layer0_outputs(9998));
    layer1_outputs(5139) <= (layer0_outputs(5068)) xor (layer0_outputs(6590));
    layer1_outputs(5140) <= '0';
    layer1_outputs(5141) <= not(layer0_outputs(7290));
    layer1_outputs(5142) <= not(layer0_outputs(9297));
    layer1_outputs(5143) <= layer0_outputs(863);
    layer1_outputs(5144) <= (layer0_outputs(2225)) or (layer0_outputs(6373));
    layer1_outputs(5145) <= layer0_outputs(5795);
    layer1_outputs(5146) <= not(layer0_outputs(9821));
    layer1_outputs(5147) <= (layer0_outputs(2004)) and not (layer0_outputs(9731));
    layer1_outputs(5148) <= not(layer0_outputs(4129));
    layer1_outputs(5149) <= layer0_outputs(1456);
    layer1_outputs(5150) <= not(layer0_outputs(6929));
    layer1_outputs(5151) <= (layer0_outputs(5812)) and (layer0_outputs(4480));
    layer1_outputs(5152) <= layer0_outputs(5048);
    layer1_outputs(5153) <= not((layer0_outputs(3864)) or (layer0_outputs(631)));
    layer1_outputs(5154) <= not((layer0_outputs(9705)) or (layer0_outputs(7736)));
    layer1_outputs(5155) <= not(layer0_outputs(400));
    layer1_outputs(5156) <= not(layer0_outputs(403)) or (layer0_outputs(9311));
    layer1_outputs(5157) <= not((layer0_outputs(7971)) xor (layer0_outputs(382)));
    layer1_outputs(5158) <= not(layer0_outputs(623));
    layer1_outputs(5159) <= not((layer0_outputs(1908)) and (layer0_outputs(7486)));
    layer1_outputs(5160) <= layer0_outputs(862);
    layer1_outputs(5161) <= layer0_outputs(9835);
    layer1_outputs(5162) <= not(layer0_outputs(2918));
    layer1_outputs(5163) <= layer0_outputs(5018);
    layer1_outputs(5164) <= (layer0_outputs(2175)) and not (layer0_outputs(1369));
    layer1_outputs(5165) <= not(layer0_outputs(2200)) or (layer0_outputs(8273));
    layer1_outputs(5166) <= '1';
    layer1_outputs(5167) <= (layer0_outputs(5722)) and not (layer0_outputs(2480));
    layer1_outputs(5168) <= (layer0_outputs(3481)) and not (layer0_outputs(4362));
    layer1_outputs(5169) <= layer0_outputs(3734);
    layer1_outputs(5170) <= not((layer0_outputs(134)) and (layer0_outputs(1476)));
    layer1_outputs(5171) <= not(layer0_outputs(9942)) or (layer0_outputs(3005));
    layer1_outputs(5172) <= not((layer0_outputs(6628)) and (layer0_outputs(2883)));
    layer1_outputs(5173) <= (layer0_outputs(3802)) and not (layer0_outputs(6295));
    layer1_outputs(5174) <= layer0_outputs(6533);
    layer1_outputs(5175) <= layer0_outputs(6964);
    layer1_outputs(5176) <= layer0_outputs(9501);
    layer1_outputs(5177) <= layer0_outputs(3656);
    layer1_outputs(5178) <= not((layer0_outputs(6855)) and (layer0_outputs(9137)));
    layer1_outputs(5179) <= not((layer0_outputs(1490)) xor (layer0_outputs(3548)));
    layer1_outputs(5180) <= (layer0_outputs(9954)) and not (layer0_outputs(8858));
    layer1_outputs(5181) <= layer0_outputs(9798);
    layer1_outputs(5182) <= not((layer0_outputs(8472)) and (layer0_outputs(3355)));
    layer1_outputs(5183) <= layer0_outputs(5600);
    layer1_outputs(5184) <= (layer0_outputs(1897)) and not (layer0_outputs(5669));
    layer1_outputs(5185) <= not(layer0_outputs(7480));
    layer1_outputs(5186) <= layer0_outputs(2064);
    layer1_outputs(5187) <= (layer0_outputs(5540)) and not (layer0_outputs(5085));
    layer1_outputs(5188) <= (layer0_outputs(9982)) and not (layer0_outputs(149));
    layer1_outputs(5189) <= not(layer0_outputs(5998));
    layer1_outputs(5190) <= (layer0_outputs(3488)) or (layer0_outputs(1035));
    layer1_outputs(5191) <= not((layer0_outputs(1403)) or (layer0_outputs(1108)));
    layer1_outputs(5192) <= layer0_outputs(7649);
    layer1_outputs(5193) <= (layer0_outputs(5539)) and not (layer0_outputs(1654));
    layer1_outputs(5194) <= '0';
    layer1_outputs(5195) <= not((layer0_outputs(7708)) or (layer0_outputs(5047)));
    layer1_outputs(5196) <= layer0_outputs(3439);
    layer1_outputs(5197) <= not(layer0_outputs(2851));
    layer1_outputs(5198) <= (layer0_outputs(7613)) and (layer0_outputs(1633));
    layer1_outputs(5199) <= not(layer0_outputs(9));
    layer1_outputs(5200) <= not(layer0_outputs(1349));
    layer1_outputs(5201) <= not(layer0_outputs(4408));
    layer1_outputs(5202) <= (layer0_outputs(5996)) and (layer0_outputs(6886));
    layer1_outputs(5203) <= (layer0_outputs(8716)) and not (layer0_outputs(2028));
    layer1_outputs(5204) <= (layer0_outputs(2672)) xor (layer0_outputs(4833));
    layer1_outputs(5205) <= (layer0_outputs(4035)) xor (layer0_outputs(1088));
    layer1_outputs(5206) <= (layer0_outputs(326)) and (layer0_outputs(1835));
    layer1_outputs(5207) <= (layer0_outputs(943)) and (layer0_outputs(6432));
    layer1_outputs(5208) <= not(layer0_outputs(8693));
    layer1_outputs(5209) <= layer0_outputs(356);
    layer1_outputs(5210) <= not(layer0_outputs(7231));
    layer1_outputs(5211) <= layer0_outputs(4125);
    layer1_outputs(5212) <= (layer0_outputs(87)) xor (layer0_outputs(3925));
    layer1_outputs(5213) <= not(layer0_outputs(242)) or (layer0_outputs(320));
    layer1_outputs(5214) <= layer0_outputs(9467);
    layer1_outputs(5215) <= not(layer0_outputs(4360)) or (layer0_outputs(1669));
    layer1_outputs(5216) <= not(layer0_outputs(6891));
    layer1_outputs(5217) <= (layer0_outputs(4509)) xor (layer0_outputs(1857));
    layer1_outputs(5218) <= not(layer0_outputs(4411)) or (layer0_outputs(6877));
    layer1_outputs(5219) <= (layer0_outputs(1533)) or (layer0_outputs(3290));
    layer1_outputs(5220) <= (layer0_outputs(7089)) or (layer0_outputs(10214));
    layer1_outputs(5221) <= not(layer0_outputs(8592));
    layer1_outputs(5222) <= not(layer0_outputs(4494));
    layer1_outputs(5223) <= layer0_outputs(1707);
    layer1_outputs(5224) <= layer0_outputs(3896);
    layer1_outputs(5225) <= (layer0_outputs(9550)) and not (layer0_outputs(1394));
    layer1_outputs(5226) <= (layer0_outputs(5730)) and (layer0_outputs(4));
    layer1_outputs(5227) <= not(layer0_outputs(8964)) or (layer0_outputs(5908));
    layer1_outputs(5228) <= not(layer0_outputs(3198));
    layer1_outputs(5229) <= (layer0_outputs(5304)) or (layer0_outputs(2563));
    layer1_outputs(5230) <= not(layer0_outputs(5156)) or (layer0_outputs(8413));
    layer1_outputs(5231) <= (layer0_outputs(1867)) and not (layer0_outputs(9689));
    layer1_outputs(5232) <= not(layer0_outputs(3902));
    layer1_outputs(5233) <= (layer0_outputs(1182)) and not (layer0_outputs(177));
    layer1_outputs(5234) <= (layer0_outputs(6604)) and not (layer0_outputs(4772));
    layer1_outputs(5235) <= (layer0_outputs(3901)) or (layer0_outputs(3792));
    layer1_outputs(5236) <= not((layer0_outputs(7235)) and (layer0_outputs(2229)));
    layer1_outputs(5237) <= not(layer0_outputs(7413)) or (layer0_outputs(6972));
    layer1_outputs(5238) <= not(layer0_outputs(5224)) or (layer0_outputs(9652));
    layer1_outputs(5239) <= not((layer0_outputs(2778)) or (layer0_outputs(5922)));
    layer1_outputs(5240) <= not(layer0_outputs(4839)) or (layer0_outputs(3350));
    layer1_outputs(5241) <= not(layer0_outputs(836)) or (layer0_outputs(5344));
    layer1_outputs(5242) <= not(layer0_outputs(9427));
    layer1_outputs(5243) <= not((layer0_outputs(6070)) or (layer0_outputs(8182)));
    layer1_outputs(5244) <= layer0_outputs(968);
    layer1_outputs(5245) <= layer0_outputs(4575);
    layer1_outputs(5246) <= (layer0_outputs(2916)) and (layer0_outputs(322));
    layer1_outputs(5247) <= layer0_outputs(1016);
    layer1_outputs(5248) <= (layer0_outputs(2569)) and (layer0_outputs(2191));
    layer1_outputs(5249) <= (layer0_outputs(8593)) and not (layer0_outputs(4584));
    layer1_outputs(5250) <= not(layer0_outputs(9581)) or (layer0_outputs(9561));
    layer1_outputs(5251) <= not(layer0_outputs(3580)) or (layer0_outputs(8337));
    layer1_outputs(5252) <= (layer0_outputs(1613)) and not (layer0_outputs(8604));
    layer1_outputs(5253) <= layer0_outputs(3254);
    layer1_outputs(5254) <= not(layer0_outputs(5936));
    layer1_outputs(5255) <= (layer0_outputs(6971)) xor (layer0_outputs(8485));
    layer1_outputs(5256) <= not((layer0_outputs(6965)) and (layer0_outputs(5918)));
    layer1_outputs(5257) <= (layer0_outputs(7714)) or (layer0_outputs(4516));
    layer1_outputs(5258) <= not(layer0_outputs(3876)) or (layer0_outputs(3776));
    layer1_outputs(5259) <= not((layer0_outputs(985)) and (layer0_outputs(8117)));
    layer1_outputs(5260) <= (layer0_outputs(9990)) and (layer0_outputs(5002));
    layer1_outputs(5261) <= (layer0_outputs(3112)) or (layer0_outputs(7576));
    layer1_outputs(5262) <= not((layer0_outputs(6642)) and (layer0_outputs(1818)));
    layer1_outputs(5263) <= not(layer0_outputs(3682));
    layer1_outputs(5264) <= not(layer0_outputs(122));
    layer1_outputs(5265) <= (layer0_outputs(6478)) and not (layer0_outputs(9276));
    layer1_outputs(5266) <= not(layer0_outputs(2640)) or (layer0_outputs(1527));
    layer1_outputs(5267) <= not((layer0_outputs(637)) and (layer0_outputs(5040)));
    layer1_outputs(5268) <= not(layer0_outputs(6120));
    layer1_outputs(5269) <= (layer0_outputs(5687)) and (layer0_outputs(6435));
    layer1_outputs(5270) <= not((layer0_outputs(6836)) xor (layer0_outputs(8562)));
    layer1_outputs(5271) <= '1';
    layer1_outputs(5272) <= (layer0_outputs(4810)) or (layer0_outputs(7108));
    layer1_outputs(5273) <= (layer0_outputs(5185)) and not (layer0_outputs(331));
    layer1_outputs(5274) <= layer0_outputs(5288);
    layer1_outputs(5275) <= not((layer0_outputs(4663)) or (layer0_outputs(6770)));
    layer1_outputs(5276) <= '0';
    layer1_outputs(5277) <= not(layer0_outputs(6434));
    layer1_outputs(5278) <= not(layer0_outputs(8388));
    layer1_outputs(5279) <= (layer0_outputs(6446)) xor (layer0_outputs(2784));
    layer1_outputs(5280) <= not(layer0_outputs(2398));
    layer1_outputs(5281) <= not(layer0_outputs(7267)) or (layer0_outputs(4342));
    layer1_outputs(5282) <= (layer0_outputs(8548)) or (layer0_outputs(1056));
    layer1_outputs(5283) <= layer0_outputs(10054);
    layer1_outputs(5284) <= (layer0_outputs(6210)) and not (layer0_outputs(10170));
    layer1_outputs(5285) <= layer0_outputs(7425);
    layer1_outputs(5286) <= not((layer0_outputs(10078)) and (layer0_outputs(5283)));
    layer1_outputs(5287) <= layer0_outputs(9665);
    layer1_outputs(5288) <= not((layer0_outputs(4305)) xor (layer0_outputs(6992)));
    layer1_outputs(5289) <= not((layer0_outputs(4878)) and (layer0_outputs(3789)));
    layer1_outputs(5290) <= not(layer0_outputs(8664));
    layer1_outputs(5291) <= not((layer0_outputs(4142)) xor (layer0_outputs(8487)));
    layer1_outputs(5292) <= (layer0_outputs(9971)) and (layer0_outputs(3991));
    layer1_outputs(5293) <= not((layer0_outputs(7180)) and (layer0_outputs(1686)));
    layer1_outputs(5294) <= not((layer0_outputs(5457)) or (layer0_outputs(101)));
    layer1_outputs(5295) <= not((layer0_outputs(9270)) or (layer0_outputs(388)));
    layer1_outputs(5296) <= not((layer0_outputs(438)) and (layer0_outputs(9638)));
    layer1_outputs(5297) <= (layer0_outputs(5145)) or (layer0_outputs(7263));
    layer1_outputs(5298) <= layer0_outputs(2675);
    layer1_outputs(5299) <= layer0_outputs(4181);
    layer1_outputs(5300) <= layer0_outputs(2043);
    layer1_outputs(5301) <= not(layer0_outputs(10076));
    layer1_outputs(5302) <= not((layer0_outputs(7518)) and (layer0_outputs(2683)));
    layer1_outputs(5303) <= not(layer0_outputs(4761));
    layer1_outputs(5304) <= (layer0_outputs(4213)) and (layer0_outputs(3521));
    layer1_outputs(5305) <= not(layer0_outputs(61));
    layer1_outputs(5306) <= (layer0_outputs(1995)) and not (layer0_outputs(5871));
    layer1_outputs(5307) <= '1';
    layer1_outputs(5308) <= '1';
    layer1_outputs(5309) <= (layer0_outputs(7624)) or (layer0_outputs(8499));
    layer1_outputs(5310) <= '1';
    layer1_outputs(5311) <= (layer0_outputs(336)) and not (layer0_outputs(695));
    layer1_outputs(5312) <= (layer0_outputs(9867)) and (layer0_outputs(3092));
    layer1_outputs(5313) <= (layer0_outputs(1363)) xor (layer0_outputs(3682));
    layer1_outputs(5314) <= not(layer0_outputs(2211));
    layer1_outputs(5315) <= not(layer0_outputs(4946)) or (layer0_outputs(4908));
    layer1_outputs(5316) <= layer0_outputs(5776);
    layer1_outputs(5317) <= not(layer0_outputs(3894));
    layer1_outputs(5318) <= (layer0_outputs(7551)) xor (layer0_outputs(5937));
    layer1_outputs(5319) <= not(layer0_outputs(8873));
    layer1_outputs(5320) <= not((layer0_outputs(7204)) xor (layer0_outputs(2205)));
    layer1_outputs(5321) <= layer0_outputs(7152);
    layer1_outputs(5322) <= layer0_outputs(1152);
    layer1_outputs(5323) <= (layer0_outputs(4965)) and (layer0_outputs(3589));
    layer1_outputs(5324) <= (layer0_outputs(3738)) and not (layer0_outputs(2066));
    layer1_outputs(5325) <= not((layer0_outputs(6223)) xor (layer0_outputs(2590)));
    layer1_outputs(5326) <= not(layer0_outputs(3857));
    layer1_outputs(5327) <= not(layer0_outputs(598)) or (layer0_outputs(103));
    layer1_outputs(5328) <= not(layer0_outputs(8272)) or (layer0_outputs(9696));
    layer1_outputs(5329) <= not(layer0_outputs(5246)) or (layer0_outputs(103));
    layer1_outputs(5330) <= not(layer0_outputs(4310));
    layer1_outputs(5331) <= not((layer0_outputs(882)) xor (layer0_outputs(7339)));
    layer1_outputs(5332) <= (layer0_outputs(6286)) and (layer0_outputs(5812));
    layer1_outputs(5333) <= not((layer0_outputs(5412)) xor (layer0_outputs(7685)));
    layer1_outputs(5334) <= layer0_outputs(7987);
    layer1_outputs(5335) <= layer0_outputs(8422);
    layer1_outputs(5336) <= not((layer0_outputs(3445)) or (layer0_outputs(1622)));
    layer1_outputs(5337) <= not(layer0_outputs(7639)) or (layer0_outputs(1332));
    layer1_outputs(5338) <= layer0_outputs(491);
    layer1_outputs(5339) <= not(layer0_outputs(10004));
    layer1_outputs(5340) <= layer0_outputs(4685);
    layer1_outputs(5341) <= not(layer0_outputs(9362)) or (layer0_outputs(3113));
    layer1_outputs(5342) <= (layer0_outputs(8240)) or (layer0_outputs(9306));
    layer1_outputs(5343) <= not((layer0_outputs(7181)) xor (layer0_outputs(4009)));
    layer1_outputs(5344) <= layer0_outputs(8649);
    layer1_outputs(5345) <= not((layer0_outputs(9050)) and (layer0_outputs(7861)));
    layer1_outputs(5346) <= '0';
    layer1_outputs(5347) <= not(layer0_outputs(2294));
    layer1_outputs(5348) <= not(layer0_outputs(6086)) or (layer0_outputs(2017));
    layer1_outputs(5349) <= not(layer0_outputs(5701)) or (layer0_outputs(2466));
    layer1_outputs(5350) <= (layer0_outputs(1298)) and not (layer0_outputs(3153));
    layer1_outputs(5351) <= not(layer0_outputs(8356)) or (layer0_outputs(3962));
    layer1_outputs(5352) <= not(layer0_outputs(7047)) or (layer0_outputs(9847));
    layer1_outputs(5353) <= not(layer0_outputs(7752));
    layer1_outputs(5354) <= not(layer0_outputs(7240));
    layer1_outputs(5355) <= not((layer0_outputs(7945)) xor (layer0_outputs(8934)));
    layer1_outputs(5356) <= layer0_outputs(8155);
    layer1_outputs(5357) <= layer0_outputs(9583);
    layer1_outputs(5358) <= '1';
    layer1_outputs(5359) <= (layer0_outputs(8557)) and not (layer0_outputs(6676));
    layer1_outputs(5360) <= layer0_outputs(9663);
    layer1_outputs(5361) <= not((layer0_outputs(303)) and (layer0_outputs(5101)));
    layer1_outputs(5362) <= '1';
    layer1_outputs(5363) <= not((layer0_outputs(8962)) and (layer0_outputs(8776)));
    layer1_outputs(5364) <= not(layer0_outputs(7063));
    layer1_outputs(5365) <= (layer0_outputs(7322)) and not (layer0_outputs(1893));
    layer1_outputs(5366) <= not(layer0_outputs(7404)) or (layer0_outputs(2852));
    layer1_outputs(5367) <= (layer0_outputs(1886)) xor (layer0_outputs(8517));
    layer1_outputs(5368) <= '1';
    layer1_outputs(5369) <= layer0_outputs(3679);
    layer1_outputs(5370) <= (layer0_outputs(5565)) or (layer0_outputs(7010));
    layer1_outputs(5371) <= not((layer0_outputs(3948)) and (layer0_outputs(4797)));
    layer1_outputs(5372) <= (layer0_outputs(377)) and not (layer0_outputs(5830));
    layer1_outputs(5373) <= not(layer0_outputs(3940)) or (layer0_outputs(1588));
    layer1_outputs(5374) <= not((layer0_outputs(8427)) xor (layer0_outputs(5696)));
    layer1_outputs(5375) <= not(layer0_outputs(1545));
    layer1_outputs(5376) <= not((layer0_outputs(2953)) xor (layer0_outputs(4440)));
    layer1_outputs(5377) <= (layer0_outputs(3873)) and (layer0_outputs(5396));
    layer1_outputs(5378) <= layer0_outputs(6687);
    layer1_outputs(5379) <= not((layer0_outputs(8568)) and (layer0_outputs(6943)));
    layer1_outputs(5380) <= layer0_outputs(577);
    layer1_outputs(5381) <= not(layer0_outputs(3052)) or (layer0_outputs(3135));
    layer1_outputs(5382) <= not(layer0_outputs(2266)) or (layer0_outputs(1998));
    layer1_outputs(5383) <= (layer0_outputs(4252)) and (layer0_outputs(7527));
    layer1_outputs(5384) <= layer0_outputs(4473);
    layer1_outputs(5385) <= layer0_outputs(140);
    layer1_outputs(5386) <= layer0_outputs(6280);
    layer1_outputs(5387) <= not(layer0_outputs(4507));
    layer1_outputs(5388) <= (layer0_outputs(9771)) and not (layer0_outputs(7146));
    layer1_outputs(5389) <= not(layer0_outputs(2728)) or (layer0_outputs(8824));
    layer1_outputs(5390) <= (layer0_outputs(4277)) and not (layer0_outputs(6659));
    layer1_outputs(5391) <= (layer0_outputs(9943)) xor (layer0_outputs(8922));
    layer1_outputs(5392) <= (layer0_outputs(7658)) and not (layer0_outputs(4727));
    layer1_outputs(5393) <= layer0_outputs(2858);
    layer1_outputs(5394) <= (layer0_outputs(7587)) and not (layer0_outputs(8739));
    layer1_outputs(5395) <= (layer0_outputs(3233)) and not (layer0_outputs(2599));
    layer1_outputs(5396) <= not(layer0_outputs(1397)) or (layer0_outputs(9995));
    layer1_outputs(5397) <= layer0_outputs(3277);
    layer1_outputs(5398) <= not(layer0_outputs(7930));
    layer1_outputs(5399) <= not((layer0_outputs(8594)) and (layer0_outputs(3173)));
    layer1_outputs(5400) <= (layer0_outputs(793)) or (layer0_outputs(6907));
    layer1_outputs(5401) <= not((layer0_outputs(1186)) xor (layer0_outputs(4576)));
    layer1_outputs(5402) <= not(layer0_outputs(6290)) or (layer0_outputs(7676));
    layer1_outputs(5403) <= layer0_outputs(7236);
    layer1_outputs(5404) <= (layer0_outputs(5610)) and not (layer0_outputs(940));
    layer1_outputs(5405) <= not(layer0_outputs(2472));
    layer1_outputs(5406) <= layer0_outputs(1353);
    layer1_outputs(5407) <= not(layer0_outputs(754)) or (layer0_outputs(9702));
    layer1_outputs(5408) <= not((layer0_outputs(3438)) xor (layer0_outputs(4971)));
    layer1_outputs(5409) <= (layer0_outputs(5831)) xor (layer0_outputs(4156));
    layer1_outputs(5410) <= not((layer0_outputs(3553)) or (layer0_outputs(10182)));
    layer1_outputs(5411) <= (layer0_outputs(2977)) xor (layer0_outputs(9521));
    layer1_outputs(5412) <= not(layer0_outputs(816));
    layer1_outputs(5413) <= not(layer0_outputs(5530));
    layer1_outputs(5414) <= not((layer0_outputs(5436)) or (layer0_outputs(1137)));
    layer1_outputs(5415) <= not(layer0_outputs(4356));
    layer1_outputs(5416) <= not((layer0_outputs(6162)) xor (layer0_outputs(7504)));
    layer1_outputs(5417) <= '1';
    layer1_outputs(5418) <= not((layer0_outputs(2680)) or (layer0_outputs(1435)));
    layer1_outputs(5419) <= not((layer0_outputs(9655)) or (layer0_outputs(3356)));
    layer1_outputs(5420) <= (layer0_outputs(8575)) and (layer0_outputs(7170));
    layer1_outputs(5421) <= not(layer0_outputs(7792));
    layer1_outputs(5422) <= layer0_outputs(5849);
    layer1_outputs(5423) <= not((layer0_outputs(299)) xor (layer0_outputs(7566)));
    layer1_outputs(5424) <= (layer0_outputs(3554)) or (layer0_outputs(2275));
    layer1_outputs(5425) <= not(layer0_outputs(4525));
    layer1_outputs(5426) <= not(layer0_outputs(10066));
    layer1_outputs(5427) <= layer0_outputs(3519);
    layer1_outputs(5428) <= layer0_outputs(4550);
    layer1_outputs(5429) <= not(layer0_outputs(6621));
    layer1_outputs(5430) <= layer0_outputs(7660);
    layer1_outputs(5431) <= (layer0_outputs(7052)) and not (layer0_outputs(1853));
    layer1_outputs(5432) <= not((layer0_outputs(4081)) or (layer0_outputs(2798)));
    layer1_outputs(5433) <= not(layer0_outputs(4414)) or (layer0_outputs(4918));
    layer1_outputs(5434) <= (layer0_outputs(1385)) xor (layer0_outputs(3201));
    layer1_outputs(5435) <= (layer0_outputs(4579)) and (layer0_outputs(601));
    layer1_outputs(5436) <= not(layer0_outputs(3056));
    layer1_outputs(5437) <= layer0_outputs(5766);
    layer1_outputs(5438) <= (layer0_outputs(1540)) or (layer0_outputs(5848));
    layer1_outputs(5439) <= not(layer0_outputs(8034)) or (layer0_outputs(9396));
    layer1_outputs(5440) <= layer0_outputs(1772);
    layer1_outputs(5441) <= not(layer0_outputs(5409));
    layer1_outputs(5442) <= not(layer0_outputs(5758));
    layer1_outputs(5443) <= not((layer0_outputs(3250)) and (layer0_outputs(2742)));
    layer1_outputs(5444) <= (layer0_outputs(4821)) or (layer0_outputs(6520));
    layer1_outputs(5445) <= not((layer0_outputs(9614)) or (layer0_outputs(6660)));
    layer1_outputs(5446) <= (layer0_outputs(5225)) and not (layer0_outputs(5166));
    layer1_outputs(5447) <= not(layer0_outputs(8433));
    layer1_outputs(5448) <= (layer0_outputs(4609)) and (layer0_outputs(8914));
    layer1_outputs(5449) <= not(layer0_outputs(7226));
    layer1_outputs(5450) <= not(layer0_outputs(5632)) or (layer0_outputs(8201));
    layer1_outputs(5451) <= not(layer0_outputs(5748));
    layer1_outputs(5452) <= (layer0_outputs(3969)) or (layer0_outputs(7939));
    layer1_outputs(5453) <= not((layer0_outputs(1832)) or (layer0_outputs(130)));
    layer1_outputs(5454) <= not(layer0_outputs(2011)) or (layer0_outputs(2846));
    layer1_outputs(5455) <= layer0_outputs(5250);
    layer1_outputs(5456) <= not(layer0_outputs(7497)) or (layer0_outputs(2084));
    layer1_outputs(5457) <= (layer0_outputs(3820)) and not (layer0_outputs(5664));
    layer1_outputs(5458) <= layer0_outputs(6371);
    layer1_outputs(5459) <= not((layer0_outputs(6763)) or (layer0_outputs(2545)));
    layer1_outputs(5460) <= layer0_outputs(9511);
    layer1_outputs(5461) <= not(layer0_outputs(7901)) or (layer0_outputs(5898));
    layer1_outputs(5462) <= layer0_outputs(4790);
    layer1_outputs(5463) <= not(layer0_outputs(3258));
    layer1_outputs(5464) <= not(layer0_outputs(5189));
    layer1_outputs(5465) <= not((layer0_outputs(811)) and (layer0_outputs(6067)));
    layer1_outputs(5466) <= layer0_outputs(4632);
    layer1_outputs(5467) <= not(layer0_outputs(5265));
    layer1_outputs(5468) <= layer0_outputs(810);
    layer1_outputs(5469) <= not(layer0_outputs(3311)) or (layer0_outputs(9911));
    layer1_outputs(5470) <= not(layer0_outputs(8727));
    layer1_outputs(5471) <= (layer0_outputs(8369)) and not (layer0_outputs(1187));
    layer1_outputs(5472) <= not((layer0_outputs(8000)) or (layer0_outputs(5613)));
    layer1_outputs(5473) <= layer0_outputs(1157);
    layer1_outputs(5474) <= (layer0_outputs(8738)) and not (layer0_outputs(6104));
    layer1_outputs(5475) <= not(layer0_outputs(8075)) or (layer0_outputs(6612));
    layer1_outputs(5476) <= not(layer0_outputs(4911));
    layer1_outputs(5477) <= layer0_outputs(5561);
    layer1_outputs(5478) <= not((layer0_outputs(3492)) and (layer0_outputs(8210)));
    layer1_outputs(5479) <= (layer0_outputs(2062)) or (layer0_outputs(183));
    layer1_outputs(5480) <= not(layer0_outputs(670));
    layer1_outputs(5481) <= not((layer0_outputs(1202)) and (layer0_outputs(9166)));
    layer1_outputs(5482) <= layer0_outputs(6025);
    layer1_outputs(5483) <= layer0_outputs(2699);
    layer1_outputs(5484) <= (layer0_outputs(711)) and (layer0_outputs(5279));
    layer1_outputs(5485) <= layer0_outputs(7719);
    layer1_outputs(5486) <= not(layer0_outputs(8622));
    layer1_outputs(5487) <= (layer0_outputs(1162)) or (layer0_outputs(7551));
    layer1_outputs(5488) <= layer0_outputs(8151);
    layer1_outputs(5489) <= layer0_outputs(9045);
    layer1_outputs(5490) <= not(layer0_outputs(2823));
    layer1_outputs(5491) <= not((layer0_outputs(8402)) or (layer0_outputs(2767)));
    layer1_outputs(5492) <= (layer0_outputs(3184)) and not (layer0_outputs(3478));
    layer1_outputs(5493) <= layer0_outputs(473);
    layer1_outputs(5494) <= not(layer0_outputs(308)) or (layer0_outputs(9795));
    layer1_outputs(5495) <= not(layer0_outputs(8592));
    layer1_outputs(5496) <= layer0_outputs(478);
    layer1_outputs(5497) <= (layer0_outputs(1746)) and not (layer0_outputs(5806));
    layer1_outputs(5498) <= not((layer0_outputs(2735)) or (layer0_outputs(4086)));
    layer1_outputs(5499) <= not(layer0_outputs(8479)) or (layer0_outputs(2587));
    layer1_outputs(5500) <= not((layer0_outputs(7072)) xor (layer0_outputs(5906)));
    layer1_outputs(5501) <= not((layer0_outputs(2297)) xor (layer0_outputs(2927)));
    layer1_outputs(5502) <= not(layer0_outputs(5264));
    layer1_outputs(5503) <= (layer0_outputs(5095)) and not (layer0_outputs(4925));
    layer1_outputs(5504) <= layer0_outputs(1886);
    layer1_outputs(5505) <= not(layer0_outputs(6029)) or (layer0_outputs(730));
    layer1_outputs(5506) <= (layer0_outputs(5051)) xor (layer0_outputs(2256));
    layer1_outputs(5507) <= (layer0_outputs(3114)) and not (layer0_outputs(1766));
    layer1_outputs(5508) <= not(layer0_outputs(8900));
    layer1_outputs(5509) <= not(layer0_outputs(813));
    layer1_outputs(5510) <= not(layer0_outputs(3471)) or (layer0_outputs(1688));
    layer1_outputs(5511) <= layer0_outputs(7459);
    layer1_outputs(5512) <= not(layer0_outputs(2237)) or (layer0_outputs(4422));
    layer1_outputs(5513) <= not((layer0_outputs(3599)) or (layer0_outputs(5011)));
    layer1_outputs(5514) <= not((layer0_outputs(9602)) xor (layer0_outputs(2468)));
    layer1_outputs(5515) <= '1';
    layer1_outputs(5516) <= (layer0_outputs(789)) and not (layer0_outputs(1913));
    layer1_outputs(5517) <= not(layer0_outputs(10207)) or (layer0_outputs(4727));
    layer1_outputs(5518) <= (layer0_outputs(9079)) and not (layer0_outputs(9672));
    layer1_outputs(5519) <= not(layer0_outputs(7483));
    layer1_outputs(5520) <= not(layer0_outputs(8018));
    layer1_outputs(5521) <= layer0_outputs(228);
    layer1_outputs(5522) <= not((layer0_outputs(6940)) xor (layer0_outputs(980)));
    layer1_outputs(5523) <= layer0_outputs(230);
    layer1_outputs(5524) <= not(layer0_outputs(542));
    layer1_outputs(5525) <= '0';
    layer1_outputs(5526) <= layer0_outputs(10143);
    layer1_outputs(5527) <= not(layer0_outputs(7398));
    layer1_outputs(5528) <= (layer0_outputs(7042)) and (layer0_outputs(3582));
    layer1_outputs(5529) <= not(layer0_outputs(9920));
    layer1_outputs(5530) <= not(layer0_outputs(8470)) or (layer0_outputs(5435));
    layer1_outputs(5531) <= layer0_outputs(7612);
    layer1_outputs(5532) <= not(layer0_outputs(9097)) or (layer0_outputs(5425));
    layer1_outputs(5533) <= (layer0_outputs(2873)) and (layer0_outputs(4686));
    layer1_outputs(5534) <= not(layer0_outputs(549));
    layer1_outputs(5535) <= layer0_outputs(8208);
    layer1_outputs(5536) <= not(layer0_outputs(3545)) or (layer0_outputs(4568));
    layer1_outputs(5537) <= not(layer0_outputs(2177)) or (layer0_outputs(8082));
    layer1_outputs(5538) <= not(layer0_outputs(6460)) or (layer0_outputs(6700));
    layer1_outputs(5539) <= (layer0_outputs(5272)) or (layer0_outputs(2639));
    layer1_outputs(5540) <= not((layer0_outputs(7103)) xor (layer0_outputs(8416)));
    layer1_outputs(5541) <= not((layer0_outputs(8870)) and (layer0_outputs(6534)));
    layer1_outputs(5542) <= (layer0_outputs(6920)) or (layer0_outputs(1537));
    layer1_outputs(5543) <= layer0_outputs(919);
    layer1_outputs(5544) <= (layer0_outputs(7681)) and not (layer0_outputs(389));
    layer1_outputs(5545) <= layer0_outputs(10113);
    layer1_outputs(5546) <= '0';
    layer1_outputs(5547) <= not((layer0_outputs(3665)) and (layer0_outputs(6878)));
    layer1_outputs(5548) <= (layer0_outputs(8902)) and (layer0_outputs(432));
    layer1_outputs(5549) <= (layer0_outputs(9281)) and not (layer0_outputs(6695));
    layer1_outputs(5550) <= not(layer0_outputs(134)) or (layer0_outputs(6317));
    layer1_outputs(5551) <= not(layer0_outputs(8860));
    layer1_outputs(5552) <= (layer0_outputs(6934)) and not (layer0_outputs(6412));
    layer1_outputs(5553) <= layer0_outputs(2149);
    layer1_outputs(5554) <= not(layer0_outputs(6933)) or (layer0_outputs(6945));
    layer1_outputs(5555) <= (layer0_outputs(5618)) and not (layer0_outputs(9851));
    layer1_outputs(5556) <= (layer0_outputs(256)) and (layer0_outputs(2416));
    layer1_outputs(5557) <= not(layer0_outputs(4109));
    layer1_outputs(5558) <= not(layer0_outputs(2784)) or (layer0_outputs(3888));
    layer1_outputs(5559) <= layer0_outputs(4015);
    layer1_outputs(5560) <= layer0_outputs(9246);
    layer1_outputs(5561) <= not(layer0_outputs(6897));
    layer1_outputs(5562) <= (layer0_outputs(110)) or (layer0_outputs(8144));
    layer1_outputs(5563) <= (layer0_outputs(5856)) and not (layer0_outputs(2582));
    layer1_outputs(5564) <= not(layer0_outputs(3523));
    layer1_outputs(5565) <= layer0_outputs(4444);
    layer1_outputs(5566) <= (layer0_outputs(9957)) xor (layer0_outputs(8446));
    layer1_outputs(5567) <= (layer0_outputs(7420)) and not (layer0_outputs(3673));
    layer1_outputs(5568) <= layer0_outputs(1143);
    layer1_outputs(5569) <= (layer0_outputs(2135)) and not (layer0_outputs(5756));
    layer1_outputs(5570) <= not(layer0_outputs(3586));
    layer1_outputs(5571) <= (layer0_outputs(8289)) xor (layer0_outputs(909));
    layer1_outputs(5572) <= (layer0_outputs(5440)) and (layer0_outputs(6463));
    layer1_outputs(5573) <= (layer0_outputs(952)) and not (layer0_outputs(2465));
    layer1_outputs(5574) <= (layer0_outputs(1070)) or (layer0_outputs(3680));
    layer1_outputs(5575) <= layer0_outputs(1923);
    layer1_outputs(5576) <= (layer0_outputs(3401)) or (layer0_outputs(3938));
    layer1_outputs(5577) <= not(layer0_outputs(9159)) or (layer0_outputs(9067));
    layer1_outputs(5578) <= not(layer0_outputs(5864)) or (layer0_outputs(5641));
    layer1_outputs(5579) <= '0';
    layer1_outputs(5580) <= (layer0_outputs(531)) xor (layer0_outputs(6416));
    layer1_outputs(5581) <= not(layer0_outputs(1896));
    layer1_outputs(5582) <= (layer0_outputs(10117)) or (layer0_outputs(8559));
    layer1_outputs(5583) <= not(layer0_outputs(8475)) or (layer0_outputs(3822));
    layer1_outputs(5584) <= not((layer0_outputs(9433)) or (layer0_outputs(1958)));
    layer1_outputs(5585) <= not(layer0_outputs(10239)) or (layer0_outputs(7807));
    layer1_outputs(5586) <= not(layer0_outputs(5541)) or (layer0_outputs(9759));
    layer1_outputs(5587) <= layer0_outputs(1821);
    layer1_outputs(5588) <= not(layer0_outputs(6908)) or (layer0_outputs(9772));
    layer1_outputs(5589) <= (layer0_outputs(9943)) and not (layer0_outputs(9641));
    layer1_outputs(5590) <= layer0_outputs(4870);
    layer1_outputs(5591) <= not((layer0_outputs(6825)) and (layer0_outputs(2808)));
    layer1_outputs(5592) <= not((layer0_outputs(2425)) or (layer0_outputs(3408)));
    layer1_outputs(5593) <= not(layer0_outputs(7479)) or (layer0_outputs(7616));
    layer1_outputs(5594) <= not(layer0_outputs(6277)) or (layer0_outputs(5042));
    layer1_outputs(5595) <= (layer0_outputs(4479)) xor (layer0_outputs(6341));
    layer1_outputs(5596) <= layer0_outputs(2442);
    layer1_outputs(5597) <= not(layer0_outputs(1646)) or (layer0_outputs(7195));
    layer1_outputs(5598) <= layer0_outputs(2372);
    layer1_outputs(5599) <= not((layer0_outputs(9840)) xor (layer0_outputs(7251)));
    layer1_outputs(5600) <= (layer0_outputs(6575)) xor (layer0_outputs(8188));
    layer1_outputs(5601) <= (layer0_outputs(3109)) xor (layer0_outputs(8630));
    layer1_outputs(5602) <= (layer0_outputs(3435)) and not (layer0_outputs(5619));
    layer1_outputs(5603) <= not(layer0_outputs(4109));
    layer1_outputs(5604) <= (layer0_outputs(2187)) and not (layer0_outputs(5611));
    layer1_outputs(5605) <= (layer0_outputs(5421)) and not (layer0_outputs(10099));
    layer1_outputs(5606) <= (layer0_outputs(9400)) xor (layer0_outputs(544));
    layer1_outputs(5607) <= (layer0_outputs(6914)) and not (layer0_outputs(2737));
    layer1_outputs(5608) <= '1';
    layer1_outputs(5609) <= (layer0_outputs(1418)) and not (layer0_outputs(6073));
    layer1_outputs(5610) <= not((layer0_outputs(708)) xor (layer0_outputs(10181)));
    layer1_outputs(5611) <= not(layer0_outputs(5887)) or (layer0_outputs(5256));
    layer1_outputs(5612) <= (layer0_outputs(2019)) and (layer0_outputs(9613));
    layer1_outputs(5613) <= layer0_outputs(9869);
    layer1_outputs(5614) <= (layer0_outputs(4897)) and not (layer0_outputs(6464));
    layer1_outputs(5615) <= not(layer0_outputs(7118)) or (layer0_outputs(8991));
    layer1_outputs(5616) <= layer0_outputs(1273);
    layer1_outputs(5617) <= (layer0_outputs(5044)) and not (layer0_outputs(6555));
    layer1_outputs(5618) <= not(layer0_outputs(7068)) or (layer0_outputs(7749));
    layer1_outputs(5619) <= not(layer0_outputs(10188));
    layer1_outputs(5620) <= (layer0_outputs(5933)) xor (layer0_outputs(2623));
    layer1_outputs(5621) <= not((layer0_outputs(3576)) xor (layer0_outputs(6665)));
    layer1_outputs(5622) <= (layer0_outputs(8962)) and (layer0_outputs(4656));
    layer1_outputs(5623) <= (layer0_outputs(2375)) or (layer0_outputs(9663));
    layer1_outputs(5624) <= not(layer0_outputs(5253)) or (layer0_outputs(2897));
    layer1_outputs(5625) <= not(layer0_outputs(4278)) or (layer0_outputs(3878));
    layer1_outputs(5626) <= (layer0_outputs(8788)) and not (layer0_outputs(9946));
    layer1_outputs(5627) <= not(layer0_outputs(6193));
    layer1_outputs(5628) <= layer0_outputs(4786);
    layer1_outputs(5629) <= layer0_outputs(4709);
    layer1_outputs(5630) <= layer0_outputs(2996);
    layer1_outputs(5631) <= (layer0_outputs(4959)) xor (layer0_outputs(9446));
    layer1_outputs(5632) <= not(layer0_outputs(6900)) or (layer0_outputs(2581));
    layer1_outputs(5633) <= (layer0_outputs(8598)) or (layer0_outputs(1982));
    layer1_outputs(5634) <= layer0_outputs(6959);
    layer1_outputs(5635) <= not(layer0_outputs(8872)) or (layer0_outputs(5518));
    layer1_outputs(5636) <= layer0_outputs(3140);
    layer1_outputs(5637) <= layer0_outputs(5017);
    layer1_outputs(5638) <= not(layer0_outputs(1967)) or (layer0_outputs(641));
    layer1_outputs(5639) <= not(layer0_outputs(2230));
    layer1_outputs(5640) <= (layer0_outputs(472)) or (layer0_outputs(204));
    layer1_outputs(5641) <= not(layer0_outputs(7842));
    layer1_outputs(5642) <= layer0_outputs(6328);
    layer1_outputs(5643) <= (layer0_outputs(6445)) and not (layer0_outputs(6125));
    layer1_outputs(5644) <= layer0_outputs(3376);
    layer1_outputs(5645) <= '1';
    layer1_outputs(5646) <= not(layer0_outputs(7753)) or (layer0_outputs(10038));
    layer1_outputs(5647) <= not(layer0_outputs(321));
    layer1_outputs(5648) <= '1';
    layer1_outputs(5649) <= layer0_outputs(8184);
    layer1_outputs(5650) <= not(layer0_outputs(8644)) or (layer0_outputs(6715));
    layer1_outputs(5651) <= not(layer0_outputs(2193)) or (layer0_outputs(4800));
    layer1_outputs(5652) <= not(layer0_outputs(9125));
    layer1_outputs(5653) <= layer0_outputs(2);
    layer1_outputs(5654) <= layer0_outputs(2898);
    layer1_outputs(5655) <= not((layer0_outputs(6396)) and (layer0_outputs(9061)));
    layer1_outputs(5656) <= layer0_outputs(9016);
    layer1_outputs(5657) <= not(layer0_outputs(172)) or (layer0_outputs(8065));
    layer1_outputs(5658) <= (layer0_outputs(8889)) or (layer0_outputs(7780));
    layer1_outputs(5659) <= (layer0_outputs(3339)) or (layer0_outputs(2624));
    layer1_outputs(5660) <= not(layer0_outputs(5860));
    layer1_outputs(5661) <= not(layer0_outputs(6459));
    layer1_outputs(5662) <= not(layer0_outputs(4023));
    layer1_outputs(5663) <= not(layer0_outputs(8299));
    layer1_outputs(5664) <= not(layer0_outputs(7950));
    layer1_outputs(5665) <= not(layer0_outputs(2000)) or (layer0_outputs(3908));
    layer1_outputs(5666) <= not(layer0_outputs(2370));
    layer1_outputs(5667) <= not((layer0_outputs(5741)) or (layer0_outputs(10167)));
    layer1_outputs(5668) <= '0';
    layer1_outputs(5669) <= not(layer0_outputs(5173));
    layer1_outputs(5670) <= not((layer0_outputs(8014)) xor (layer0_outputs(11)));
    layer1_outputs(5671) <= (layer0_outputs(537)) or (layer0_outputs(7362));
    layer1_outputs(5672) <= (layer0_outputs(4810)) xor (layer0_outputs(4620));
    layer1_outputs(5673) <= (layer0_outputs(2954)) and (layer0_outputs(3002));
    layer1_outputs(5674) <= not(layer0_outputs(7186)) or (layer0_outputs(7885));
    layer1_outputs(5675) <= (layer0_outputs(9981)) and not (layer0_outputs(7139));
    layer1_outputs(5676) <= not(layer0_outputs(455));
    layer1_outputs(5677) <= (layer0_outputs(1517)) and not (layer0_outputs(6116));
    layer1_outputs(5678) <= not(layer0_outputs(2057));
    layer1_outputs(5679) <= not(layer0_outputs(7899));
    layer1_outputs(5680) <= layer0_outputs(4488);
    layer1_outputs(5681) <= not(layer0_outputs(5527));
    layer1_outputs(5682) <= not((layer0_outputs(1538)) and (layer0_outputs(7505)));
    layer1_outputs(5683) <= not(layer0_outputs(7121));
    layer1_outputs(5684) <= (layer0_outputs(7656)) xor (layer0_outputs(8847));
    layer1_outputs(5685) <= not((layer0_outputs(5909)) or (layer0_outputs(3083)));
    layer1_outputs(5686) <= not(layer0_outputs(9174)) or (layer0_outputs(9161));
    layer1_outputs(5687) <= (layer0_outputs(2628)) and not (layer0_outputs(1952));
    layer1_outputs(5688) <= not(layer0_outputs(2012)) or (layer0_outputs(9167));
    layer1_outputs(5689) <= (layer0_outputs(4735)) and (layer0_outputs(9059));
    layer1_outputs(5690) <= not(layer0_outputs(8925));
    layer1_outputs(5691) <= not(layer0_outputs(1288));
    layer1_outputs(5692) <= (layer0_outputs(9830)) or (layer0_outputs(2046));
    layer1_outputs(5693) <= (layer0_outputs(8466)) and not (layer0_outputs(894));
    layer1_outputs(5694) <= not(layer0_outputs(5176)) or (layer0_outputs(8356));
    layer1_outputs(5695) <= (layer0_outputs(266)) xor (layer0_outputs(6211));
    layer1_outputs(5696) <= not(layer0_outputs(3431));
    layer1_outputs(5697) <= layer0_outputs(167);
    layer1_outputs(5698) <= layer0_outputs(8340);
    layer1_outputs(5699) <= (layer0_outputs(714)) and not (layer0_outputs(4689));
    layer1_outputs(5700) <= (layer0_outputs(10119)) and not (layer0_outputs(4835));
    layer1_outputs(5701) <= not(layer0_outputs(7809));
    layer1_outputs(5702) <= not(layer0_outputs(4826));
    layer1_outputs(5703) <= (layer0_outputs(5767)) and not (layer0_outputs(137));
    layer1_outputs(5704) <= (layer0_outputs(954)) xor (layer0_outputs(5656));
    layer1_outputs(5705) <= not(layer0_outputs(5637));
    layer1_outputs(5706) <= (layer0_outputs(9793)) and not (layer0_outputs(5785));
    layer1_outputs(5707) <= (layer0_outputs(6469)) and (layer0_outputs(9332));
    layer1_outputs(5708) <= layer0_outputs(7075);
    layer1_outputs(5709) <= not(layer0_outputs(8761)) or (layer0_outputs(6723));
    layer1_outputs(5710) <= layer0_outputs(9885);
    layer1_outputs(5711) <= not((layer0_outputs(9662)) xor (layer0_outputs(1041)));
    layer1_outputs(5712) <= not(layer0_outputs(777)) or (layer0_outputs(560));
    layer1_outputs(5713) <= not((layer0_outputs(367)) and (layer0_outputs(7225)));
    layer1_outputs(5714) <= not(layer0_outputs(3698)) or (layer0_outputs(5651));
    layer1_outputs(5715) <= not(layer0_outputs(4342));
    layer1_outputs(5716) <= '1';
    layer1_outputs(5717) <= not(layer0_outputs(7890));
    layer1_outputs(5718) <= (layer0_outputs(6193)) and not (layer0_outputs(8008));
    layer1_outputs(5719) <= not((layer0_outputs(4422)) and (layer0_outputs(4776)));
    layer1_outputs(5720) <= not(layer0_outputs(2983));
    layer1_outputs(5721) <= (layer0_outputs(3209)) and (layer0_outputs(689));
    layer1_outputs(5722) <= not(layer0_outputs(2820));
    layer1_outputs(5723) <= not(layer0_outputs(4680));
    layer1_outputs(5724) <= (layer0_outputs(2289)) or (layer0_outputs(9233));
    layer1_outputs(5725) <= not(layer0_outputs(1445));
    layer1_outputs(5726) <= not(layer0_outputs(3648)) or (layer0_outputs(8376));
    layer1_outputs(5727) <= (layer0_outputs(5275)) or (layer0_outputs(9387));
    layer1_outputs(5728) <= not(layer0_outputs(6561)) or (layer0_outputs(8001));
    layer1_outputs(5729) <= not(layer0_outputs(7300)) or (layer0_outputs(9263));
    layer1_outputs(5730) <= not(layer0_outputs(4763));
    layer1_outputs(5731) <= layer0_outputs(3183);
    layer1_outputs(5732) <= not((layer0_outputs(8668)) and (layer0_outputs(2369)));
    layer1_outputs(5733) <= not(layer0_outputs(9017));
    layer1_outputs(5734) <= (layer0_outputs(4221)) and not (layer0_outputs(7841));
    layer1_outputs(5735) <= (layer0_outputs(7071)) and not (layer0_outputs(5746));
    layer1_outputs(5736) <= not((layer0_outputs(3039)) or (layer0_outputs(1174)));
    layer1_outputs(5737) <= not(layer0_outputs(6001));
    layer1_outputs(5738) <= not(layer0_outputs(6821));
    layer1_outputs(5739) <= not(layer0_outputs(1384));
    layer1_outputs(5740) <= not(layer0_outputs(9231));
    layer1_outputs(5741) <= layer0_outputs(3592);
    layer1_outputs(5742) <= not(layer0_outputs(3004));
    layer1_outputs(5743) <= layer0_outputs(1733);
    layer1_outputs(5744) <= layer0_outputs(1827);
    layer1_outputs(5745) <= not(layer0_outputs(9028)) or (layer0_outputs(737));
    layer1_outputs(5746) <= (layer0_outputs(1233)) and not (layer0_outputs(5281));
    layer1_outputs(5747) <= not((layer0_outputs(8887)) or (layer0_outputs(7006)));
    layer1_outputs(5748) <= not(layer0_outputs(4666));
    layer1_outputs(5749) <= (layer0_outputs(6154)) and (layer0_outputs(3772));
    layer1_outputs(5750) <= not(layer0_outputs(4038)) or (layer0_outputs(9791));
    layer1_outputs(5751) <= not((layer0_outputs(3755)) and (layer0_outputs(6424)));
    layer1_outputs(5752) <= '0';
    layer1_outputs(5753) <= not(layer0_outputs(3572)) or (layer0_outputs(5611));
    layer1_outputs(5754) <= (layer0_outputs(1291)) and not (layer0_outputs(4639));
    layer1_outputs(5755) <= not(layer0_outputs(7909));
    layer1_outputs(5756) <= (layer0_outputs(5187)) and not (layer0_outputs(8457));
    layer1_outputs(5757) <= layer0_outputs(1098);
    layer1_outputs(5758) <= layer0_outputs(2028);
    layer1_outputs(5759) <= (layer0_outputs(1016)) and not (layer0_outputs(8088));
    layer1_outputs(5760) <= layer0_outputs(9806);
    layer1_outputs(5761) <= not((layer0_outputs(1470)) or (layer0_outputs(7086)));
    layer1_outputs(5762) <= not(layer0_outputs(6766));
    layer1_outputs(5763) <= not((layer0_outputs(4270)) or (layer0_outputs(7437)));
    layer1_outputs(5764) <= not(layer0_outputs(5803));
    layer1_outputs(5765) <= not((layer0_outputs(2263)) and (layer0_outputs(350)));
    layer1_outputs(5766) <= (layer0_outputs(5309)) or (layer0_outputs(8269));
    layer1_outputs(5767) <= (layer0_outputs(8033)) or (layer0_outputs(5853));
    layer1_outputs(5768) <= '0';
    layer1_outputs(5769) <= not(layer0_outputs(6242)) or (layer0_outputs(7610));
    layer1_outputs(5770) <= not(layer0_outputs(8465));
    layer1_outputs(5771) <= not(layer0_outputs(8242));
    layer1_outputs(5772) <= not(layer0_outputs(2022)) or (layer0_outputs(6469));
    layer1_outputs(5773) <= (layer0_outputs(4977)) and not (layer0_outputs(9287));
    layer1_outputs(5774) <= layer0_outputs(9789);
    layer1_outputs(5775) <= (layer0_outputs(3090)) and not (layer0_outputs(1734));
    layer1_outputs(5776) <= not((layer0_outputs(6081)) xor (layer0_outputs(5780)));
    layer1_outputs(5777) <= (layer0_outputs(7275)) and not (layer0_outputs(3985));
    layer1_outputs(5778) <= (layer0_outputs(4555)) or (layer0_outputs(2013));
    layer1_outputs(5779) <= not(layer0_outputs(3260));
    layer1_outputs(5780) <= not(layer0_outputs(9868));
    layer1_outputs(5781) <= not(layer0_outputs(47)) or (layer0_outputs(525));
    layer1_outputs(5782) <= layer0_outputs(584);
    layer1_outputs(5783) <= not(layer0_outputs(1018));
    layer1_outputs(5784) <= (layer0_outputs(1734)) or (layer0_outputs(2689));
    layer1_outputs(5785) <= (layer0_outputs(9431)) and (layer0_outputs(5957));
    layer1_outputs(5786) <= not((layer0_outputs(9407)) and (layer0_outputs(9628)));
    layer1_outputs(5787) <= (layer0_outputs(8629)) and (layer0_outputs(7315));
    layer1_outputs(5788) <= not(layer0_outputs(4186));
    layer1_outputs(5789) <= layer0_outputs(8058);
    layer1_outputs(5790) <= not((layer0_outputs(1972)) or (layer0_outputs(8014)));
    layer1_outputs(5791) <= layer0_outputs(8520);
    layer1_outputs(5792) <= not(layer0_outputs(6165));
    layer1_outputs(5793) <= not((layer0_outputs(4642)) or (layer0_outputs(839)));
    layer1_outputs(5794) <= (layer0_outputs(9040)) xor (layer0_outputs(6865));
    layer1_outputs(5795) <= not((layer0_outputs(7530)) or (layer0_outputs(8754)));
    layer1_outputs(5796) <= not(layer0_outputs(3723));
    layer1_outputs(5797) <= layer0_outputs(6199);
    layer1_outputs(5798) <= not((layer0_outputs(3300)) xor (layer0_outputs(3341)));
    layer1_outputs(5799) <= (layer0_outputs(4274)) and not (layer0_outputs(8280));
    layer1_outputs(5800) <= (layer0_outputs(969)) and (layer0_outputs(234));
    layer1_outputs(5801) <= not(layer0_outputs(2533)) or (layer0_outputs(4602));
    layer1_outputs(5802) <= layer0_outputs(284);
    layer1_outputs(5803) <= (layer0_outputs(3436)) and not (layer0_outputs(379));
    layer1_outputs(5804) <= (layer0_outputs(7966)) or (layer0_outputs(3814));
    layer1_outputs(5805) <= layer0_outputs(1683);
    layer1_outputs(5806) <= not(layer0_outputs(7248)) or (layer0_outputs(61));
    layer1_outputs(5807) <= (layer0_outputs(2373)) or (layer0_outputs(10082));
    layer1_outputs(5808) <= (layer0_outputs(9400)) and not (layer0_outputs(988));
    layer1_outputs(5809) <= (layer0_outputs(3082)) and (layer0_outputs(6144));
    layer1_outputs(5810) <= (layer0_outputs(9951)) and not (layer0_outputs(6066));
    layer1_outputs(5811) <= (layer0_outputs(1350)) and (layer0_outputs(3066));
    layer1_outputs(5812) <= not((layer0_outputs(9293)) and (layer0_outputs(1158)));
    layer1_outputs(5813) <= (layer0_outputs(5289)) or (layer0_outputs(3911));
    layer1_outputs(5814) <= (layer0_outputs(779)) and not (layer0_outputs(4904));
    layer1_outputs(5815) <= layer0_outputs(2866);
    layer1_outputs(5816) <= not(layer0_outputs(10151));
    layer1_outputs(5817) <= not(layer0_outputs(7536)) or (layer0_outputs(3257));
    layer1_outputs(5818) <= not(layer0_outputs(2628));
    layer1_outputs(5819) <= not(layer0_outputs(5171));
    layer1_outputs(5820) <= (layer0_outputs(770)) and (layer0_outputs(8833));
    layer1_outputs(5821) <= (layer0_outputs(9745)) and (layer0_outputs(5077));
    layer1_outputs(5822) <= not((layer0_outputs(3196)) xor (layer0_outputs(5593)));
    layer1_outputs(5823) <= (layer0_outputs(6579)) xor (layer0_outputs(2410));
    layer1_outputs(5824) <= layer0_outputs(5241);
    layer1_outputs(5825) <= not(layer0_outputs(1625));
    layer1_outputs(5826) <= layer0_outputs(2254);
    layer1_outputs(5827) <= layer0_outputs(2962);
    layer1_outputs(5828) <= not((layer0_outputs(2577)) and (layer0_outputs(166)));
    layer1_outputs(5829) <= (layer0_outputs(5851)) and (layer0_outputs(7337));
    layer1_outputs(5830) <= (layer0_outputs(2316)) or (layer0_outputs(8486));
    layer1_outputs(5831) <= layer0_outputs(5659);
    layer1_outputs(5832) <= (layer0_outputs(9145)) xor (layer0_outputs(578));
    layer1_outputs(5833) <= not(layer0_outputs(4283));
    layer1_outputs(5834) <= layer0_outputs(7531);
    layer1_outputs(5835) <= not(layer0_outputs(4881));
    layer1_outputs(5836) <= layer0_outputs(5192);
    layer1_outputs(5837) <= not((layer0_outputs(7471)) xor (layer0_outputs(5690)));
    layer1_outputs(5838) <= not(layer0_outputs(9828)) or (layer0_outputs(8945));
    layer1_outputs(5839) <= layer0_outputs(8323);
    layer1_outputs(5840) <= '0';
    layer1_outputs(5841) <= not((layer0_outputs(1953)) xor (layer0_outputs(5542)));
    layer1_outputs(5842) <= not(layer0_outputs(2287));
    layer1_outputs(5843) <= layer0_outputs(5880);
    layer1_outputs(5844) <= layer0_outputs(9642);
    layer1_outputs(5845) <= (layer0_outputs(4388)) and not (layer0_outputs(6007));
    layer1_outputs(5846) <= not(layer0_outputs(726));
    layer1_outputs(5847) <= layer0_outputs(8363);
    layer1_outputs(5848) <= (layer0_outputs(9059)) and not (layer0_outputs(4172));
    layer1_outputs(5849) <= (layer0_outputs(2724)) or (layer0_outputs(2369));
    layer1_outputs(5850) <= not((layer0_outputs(4613)) or (layer0_outputs(848)));
    layer1_outputs(5851) <= not(layer0_outputs(8171));
    layer1_outputs(5852) <= (layer0_outputs(8869)) or (layer0_outputs(9562));
    layer1_outputs(5853) <= (layer0_outputs(7120)) and not (layer0_outputs(1651));
    layer1_outputs(5854) <= '1';
    layer1_outputs(5855) <= not(layer0_outputs(2568)) or (layer0_outputs(7455));
    layer1_outputs(5856) <= layer0_outputs(6374);
    layer1_outputs(5857) <= (layer0_outputs(1747)) and (layer0_outputs(5215));
    layer1_outputs(5858) <= layer0_outputs(9537);
    layer1_outputs(5859) <= layer0_outputs(2559);
    layer1_outputs(5860) <= (layer0_outputs(2120)) or (layer0_outputs(6185));
    layer1_outputs(5861) <= not((layer0_outputs(7926)) and (layer0_outputs(8711)));
    layer1_outputs(5862) <= not(layer0_outputs(176)) or (layer0_outputs(6024));
    layer1_outputs(5863) <= not((layer0_outputs(7508)) xor (layer0_outputs(8499)));
    layer1_outputs(5864) <= not(layer0_outputs(2608));
    layer1_outputs(5865) <= (layer0_outputs(9637)) and (layer0_outputs(4561));
    layer1_outputs(5866) <= not((layer0_outputs(7447)) xor (layer0_outputs(3467)));
    layer1_outputs(5867) <= '1';
    layer1_outputs(5868) <= not(layer0_outputs(9728));
    layer1_outputs(5869) <= not(layer0_outputs(7689));
    layer1_outputs(5870) <= not((layer0_outputs(4085)) or (layer0_outputs(241)));
    layer1_outputs(5871) <= (layer0_outputs(1750)) and not (layer0_outputs(2363));
    layer1_outputs(5872) <= (layer0_outputs(7635)) or (layer0_outputs(8852));
    layer1_outputs(5873) <= (layer0_outputs(3488)) and not (layer0_outputs(894));
    layer1_outputs(5874) <= (layer0_outputs(2749)) or (layer0_outputs(2319));
    layer1_outputs(5875) <= not((layer0_outputs(1987)) xor (layer0_outputs(737)));
    layer1_outputs(5876) <= (layer0_outputs(1975)) or (layer0_outputs(3229));
    layer1_outputs(5877) <= layer0_outputs(3147);
    layer1_outputs(5878) <= not(layer0_outputs(8146));
    layer1_outputs(5879) <= layer0_outputs(8997);
    layer1_outputs(5880) <= '1';
    layer1_outputs(5881) <= not((layer0_outputs(6457)) and (layer0_outputs(4221)));
    layer1_outputs(5882) <= not((layer0_outputs(8175)) and (layer0_outputs(6003)));
    layer1_outputs(5883) <= not(layer0_outputs(1875)) or (layer0_outputs(5155));
    layer1_outputs(5884) <= not((layer0_outputs(1086)) or (layer0_outputs(6984)));
    layer1_outputs(5885) <= (layer0_outputs(8200)) or (layer0_outputs(3282));
    layer1_outputs(5886) <= not((layer0_outputs(5574)) and (layer0_outputs(7027)));
    layer1_outputs(5887) <= not(layer0_outputs(3786));
    layer1_outputs(5888) <= (layer0_outputs(4443)) or (layer0_outputs(3464));
    layer1_outputs(5889) <= (layer0_outputs(6581)) or (layer0_outputs(1485));
    layer1_outputs(5890) <= layer0_outputs(5224);
    layer1_outputs(5891) <= not(layer0_outputs(1507));
    layer1_outputs(5892) <= layer0_outputs(9030);
    layer1_outputs(5893) <= not(layer0_outputs(3539));
    layer1_outputs(5894) <= not(layer0_outputs(2748));
    layer1_outputs(5895) <= not(layer0_outputs(9546));
    layer1_outputs(5896) <= not(layer0_outputs(4998));
    layer1_outputs(5897) <= not(layer0_outputs(9978));
    layer1_outputs(5898) <= (layer0_outputs(1801)) and (layer0_outputs(3688));
    layer1_outputs(5899) <= (layer0_outputs(2281)) and not (layer0_outputs(282));
    layer1_outputs(5900) <= layer0_outputs(9842);
    layer1_outputs(5901) <= (layer0_outputs(9290)) and not (layer0_outputs(5532));
    layer1_outputs(5902) <= (layer0_outputs(943)) and not (layer0_outputs(5648));
    layer1_outputs(5903) <= not(layer0_outputs(8497));
    layer1_outputs(5904) <= (layer0_outputs(106)) and not (layer0_outputs(10225));
    layer1_outputs(5905) <= layer0_outputs(2380);
    layer1_outputs(5906) <= not(layer0_outputs(196)) or (layer0_outputs(144));
    layer1_outputs(5907) <= not((layer0_outputs(518)) and (layer0_outputs(4270)));
    layer1_outputs(5908) <= layer0_outputs(9975);
    layer1_outputs(5909) <= layer0_outputs(9844);
    layer1_outputs(5910) <= not((layer0_outputs(5533)) and (layer0_outputs(5552)));
    layer1_outputs(5911) <= layer0_outputs(5536);
    layer1_outputs(5912) <= not((layer0_outputs(5275)) or (layer0_outputs(5775)));
    layer1_outputs(5913) <= not(layer0_outputs(3136)) or (layer0_outputs(7270));
    layer1_outputs(5914) <= not(layer0_outputs(6927));
    layer1_outputs(5915) <= (layer0_outputs(740)) and (layer0_outputs(9670));
    layer1_outputs(5916) <= not(layer0_outputs(2698));
    layer1_outputs(5917) <= not(layer0_outputs(10044)) or (layer0_outputs(4353));
    layer1_outputs(5918) <= '0';
    layer1_outputs(5919) <= layer0_outputs(7919);
    layer1_outputs(5920) <= not((layer0_outputs(9225)) or (layer0_outputs(1706)));
    layer1_outputs(5921) <= (layer0_outputs(8179)) xor (layer0_outputs(7648));
    layer1_outputs(5922) <= not(layer0_outputs(3060)) or (layer0_outputs(805));
    layer1_outputs(5923) <= layer0_outputs(7574);
    layer1_outputs(5924) <= (layer0_outputs(9250)) and not (layer0_outputs(6252));
    layer1_outputs(5925) <= layer0_outputs(1229);
    layer1_outputs(5926) <= not(layer0_outputs(2987)) or (layer0_outputs(728));
    layer1_outputs(5927) <= '1';
    layer1_outputs(5928) <= (layer0_outputs(9817)) or (layer0_outputs(6119));
    layer1_outputs(5929) <= (layer0_outputs(7376)) and (layer0_outputs(8488));
    layer1_outputs(5930) <= (layer0_outputs(5539)) xor (layer0_outputs(2199));
    layer1_outputs(5931) <= not(layer0_outputs(3303));
    layer1_outputs(5932) <= not((layer0_outputs(2600)) xor (layer0_outputs(330)));
    layer1_outputs(5933) <= (layer0_outputs(339)) xor (layer0_outputs(6988));
    layer1_outputs(5934) <= (layer0_outputs(10035)) and not (layer0_outputs(891));
    layer1_outputs(5935) <= (layer0_outputs(2696)) and not (layer0_outputs(3206));
    layer1_outputs(5936) <= (layer0_outputs(7691)) and not (layer0_outputs(3598));
    layer1_outputs(5937) <= not(layer0_outputs(5829));
    layer1_outputs(5938) <= not((layer0_outputs(7716)) xor (layer0_outputs(1425)));
    layer1_outputs(5939) <= layer0_outputs(4831);
    layer1_outputs(5940) <= (layer0_outputs(6431)) and (layer0_outputs(8615));
    layer1_outputs(5941) <= (layer0_outputs(6297)) and (layer0_outputs(778));
    layer1_outputs(5942) <= not(layer0_outputs(9647));
    layer1_outputs(5943) <= not(layer0_outputs(484)) or (layer0_outputs(3754));
    layer1_outputs(5944) <= layer0_outputs(11);
    layer1_outputs(5945) <= layer0_outputs(5491);
    layer1_outputs(5946) <= (layer0_outputs(3663)) and not (layer0_outputs(5491));
    layer1_outputs(5947) <= (layer0_outputs(8297)) and not (layer0_outputs(1895));
    layer1_outputs(5948) <= not(layer0_outputs(6627)) or (layer0_outputs(8372));
    layer1_outputs(5949) <= not((layer0_outputs(2809)) xor (layer0_outputs(2618)));
    layer1_outputs(5950) <= layer0_outputs(4824);
    layer1_outputs(5951) <= not(layer0_outputs(5000)) or (layer0_outputs(6393));
    layer1_outputs(5952) <= '1';
    layer1_outputs(5953) <= not(layer0_outputs(3251)) or (layer0_outputs(84));
    layer1_outputs(5954) <= layer0_outputs(6799);
    layer1_outputs(5955) <= (layer0_outputs(2149)) xor (layer0_outputs(4452));
    layer1_outputs(5956) <= layer0_outputs(6769);
    layer1_outputs(5957) <= not(layer0_outputs(9694));
    layer1_outputs(5958) <= not(layer0_outputs(4154));
    layer1_outputs(5959) <= (layer0_outputs(6134)) or (layer0_outputs(7004));
    layer1_outputs(5960) <= (layer0_outputs(7788)) and not (layer0_outputs(7080));
    layer1_outputs(5961) <= (layer0_outputs(6857)) xor (layer0_outputs(1048));
    layer1_outputs(5962) <= not((layer0_outputs(9715)) and (layer0_outputs(876)));
    layer1_outputs(5963) <= not(layer0_outputs(7355));
    layer1_outputs(5964) <= not(layer0_outputs(476)) or (layer0_outputs(5714));
    layer1_outputs(5965) <= not((layer0_outputs(2836)) xor (layer0_outputs(3404)));
    layer1_outputs(5966) <= (layer0_outputs(2634)) and not (layer0_outputs(2907));
    layer1_outputs(5967) <= not(layer0_outputs(4672));
    layer1_outputs(5968) <= layer0_outputs(7253);
    layer1_outputs(5969) <= (layer0_outputs(700)) and not (layer0_outputs(7016));
    layer1_outputs(5970) <= not(layer0_outputs(5109)) or (layer0_outputs(5822));
    layer1_outputs(5971) <= not((layer0_outputs(9952)) or (layer0_outputs(441)));
    layer1_outputs(5972) <= not(layer0_outputs(7604)) or (layer0_outputs(6501));
    layer1_outputs(5973) <= not(layer0_outputs(6593));
    layer1_outputs(5974) <= layer0_outputs(7826);
    layer1_outputs(5975) <= not((layer0_outputs(5516)) and (layer0_outputs(2532)));
    layer1_outputs(5976) <= not((layer0_outputs(5342)) xor (layer0_outputs(9284)));
    layer1_outputs(5977) <= layer0_outputs(9350);
    layer1_outputs(5978) <= not(layer0_outputs(280)) or (layer0_outputs(7671));
    layer1_outputs(5979) <= (layer0_outputs(677)) or (layer0_outputs(7396));
    layer1_outputs(5980) <= not((layer0_outputs(2151)) or (layer0_outputs(4357)));
    layer1_outputs(5981) <= not((layer0_outputs(2876)) xor (layer0_outputs(9146)));
    layer1_outputs(5982) <= (layer0_outputs(3423)) xor (layer0_outputs(2145));
    layer1_outputs(5983) <= not((layer0_outputs(9808)) or (layer0_outputs(1253)));
    layer1_outputs(5984) <= layer0_outputs(16);
    layer1_outputs(5985) <= layer0_outputs(1977);
    layer1_outputs(5986) <= (layer0_outputs(1413)) and not (layer0_outputs(9676));
    layer1_outputs(5987) <= not((layer0_outputs(8028)) or (layer0_outputs(9018)));
    layer1_outputs(5988) <= not(layer0_outputs(339));
    layer1_outputs(5989) <= not((layer0_outputs(1439)) xor (layer0_outputs(68)));
    layer1_outputs(5990) <= not(layer0_outputs(7777)) or (layer0_outputs(9073));
    layer1_outputs(5991) <= '0';
    layer1_outputs(5992) <= not(layer0_outputs(4926));
    layer1_outputs(5993) <= layer0_outputs(2725);
    layer1_outputs(5994) <= '1';
    layer1_outputs(5995) <= not(layer0_outputs(1191));
    layer1_outputs(5996) <= not((layer0_outputs(3574)) or (layer0_outputs(5496)));
    layer1_outputs(5997) <= not(layer0_outputs(8255));
    layer1_outputs(5998) <= not(layer0_outputs(1830)) or (layer0_outputs(3421));
    layer1_outputs(5999) <= not(layer0_outputs(4183));
    layer1_outputs(6000) <= not(layer0_outputs(1150)) or (layer0_outputs(2025));
    layer1_outputs(6001) <= (layer0_outputs(1967)) and not (layer0_outputs(6225));
    layer1_outputs(6002) <= not((layer0_outputs(4387)) or (layer0_outputs(9929)));
    layer1_outputs(6003) <= (layer0_outputs(4061)) and (layer0_outputs(3166));
    layer1_outputs(6004) <= not(layer0_outputs(5725)) or (layer0_outputs(6919));
    layer1_outputs(6005) <= (layer0_outputs(5970)) and (layer0_outputs(8199));
    layer1_outputs(6006) <= not((layer0_outputs(6153)) or (layer0_outputs(3537)));
    layer1_outputs(6007) <= (layer0_outputs(8401)) and (layer0_outputs(4135));
    layer1_outputs(6008) <= not(layer0_outputs(5835));
    layer1_outputs(6009) <= '1';
    layer1_outputs(6010) <= '1';
    layer1_outputs(6011) <= not(layer0_outputs(750));
    layer1_outputs(6012) <= not(layer0_outputs(1461));
    layer1_outputs(6013) <= (layer0_outputs(98)) and not (layer0_outputs(5895));
    layer1_outputs(6014) <= layer0_outputs(6934);
    layer1_outputs(6015) <= layer0_outputs(2336);
    layer1_outputs(6016) <= not((layer0_outputs(2279)) or (layer0_outputs(3856)));
    layer1_outputs(6017) <= (layer0_outputs(8714)) and not (layer0_outputs(10227));
    layer1_outputs(6018) <= (layer0_outputs(3817)) xor (layer0_outputs(4199));
    layer1_outputs(6019) <= (layer0_outputs(2805)) and not (layer0_outputs(5827));
    layer1_outputs(6020) <= not(layer0_outputs(2839));
    layer1_outputs(6021) <= not((layer0_outputs(7952)) and (layer0_outputs(5125)));
    layer1_outputs(6022) <= (layer0_outputs(9229)) and not (layer0_outputs(6691));
    layer1_outputs(6023) <= layer0_outputs(1716);
    layer1_outputs(6024) <= (layer0_outputs(3110)) or (layer0_outputs(516));
    layer1_outputs(6025) <= (layer0_outputs(7178)) and (layer0_outputs(3096));
    layer1_outputs(6026) <= (layer0_outputs(8469)) and (layer0_outputs(5460));
    layer1_outputs(6027) <= not((layer0_outputs(4702)) xor (layer0_outputs(1079)));
    layer1_outputs(6028) <= (layer0_outputs(2804)) or (layer0_outputs(9510));
    layer1_outputs(6029) <= not((layer0_outputs(4717)) and (layer0_outputs(3418)));
    layer1_outputs(6030) <= not(layer0_outputs(7477)) or (layer0_outputs(4880));
    layer1_outputs(6031) <= not(layer0_outputs(8245));
    layer1_outputs(6032) <= (layer0_outputs(6112)) and not (layer0_outputs(6013));
    layer1_outputs(6033) <= not(layer0_outputs(4180)) or (layer0_outputs(2221));
    layer1_outputs(6034) <= not(layer0_outputs(3225));
    layer1_outputs(6035) <= (layer0_outputs(484)) and (layer0_outputs(1523));
    layer1_outputs(6036) <= not(layer0_outputs(8262));
    layer1_outputs(6037) <= (layer0_outputs(8342)) xor (layer0_outputs(3363));
    layer1_outputs(6038) <= layer0_outputs(8138);
    layer1_outputs(6039) <= not(layer0_outputs(859)) or (layer0_outputs(2457));
    layer1_outputs(6040) <= layer0_outputs(6569);
    layer1_outputs(6041) <= not(layer0_outputs(1573)) or (layer0_outputs(1335));
    layer1_outputs(6042) <= (layer0_outputs(8950)) and not (layer0_outputs(7703));
    layer1_outputs(6043) <= not(layer0_outputs(1917));
    layer1_outputs(6044) <= not(layer0_outputs(5568));
    layer1_outputs(6045) <= not((layer0_outputs(7000)) and (layer0_outputs(2243)));
    layer1_outputs(6046) <= (layer0_outputs(7256)) xor (layer0_outputs(3440));
    layer1_outputs(6047) <= not(layer0_outputs(473));
    layer1_outputs(6048) <= layer0_outputs(4803);
    layer1_outputs(6049) <= not((layer0_outputs(5099)) and (layer0_outputs(6880)));
    layer1_outputs(6050) <= not(layer0_outputs(1720));
    layer1_outputs(6051) <= not((layer0_outputs(2821)) xor (layer0_outputs(7507)));
    layer1_outputs(6052) <= not(layer0_outputs(8888));
    layer1_outputs(6053) <= (layer0_outputs(8654)) or (layer0_outputs(7654));
    layer1_outputs(6054) <= not(layer0_outputs(9346));
    layer1_outputs(6055) <= (layer0_outputs(6290)) and not (layer0_outputs(6145));
    layer1_outputs(6056) <= not(layer0_outputs(6665)) or (layer0_outputs(8704));
    layer1_outputs(6057) <= not((layer0_outputs(4365)) or (layer0_outputs(1090)));
    layer1_outputs(6058) <= (layer0_outputs(2242)) and not (layer0_outputs(3703));
    layer1_outputs(6059) <= not(layer0_outputs(9436));
    layer1_outputs(6060) <= (layer0_outputs(1751)) xor (layer0_outputs(7532));
    layer1_outputs(6061) <= not(layer0_outputs(5523)) or (layer0_outputs(6117));
    layer1_outputs(6062) <= (layer0_outputs(6187)) xor (layer0_outputs(4390));
    layer1_outputs(6063) <= not(layer0_outputs(1642));
    layer1_outputs(6064) <= (layer0_outputs(3219)) or (layer0_outputs(2349));
    layer1_outputs(6065) <= (layer0_outputs(3316)) xor (layer0_outputs(2890));
    layer1_outputs(6066) <= not(layer0_outputs(502));
    layer1_outputs(6067) <= layer0_outputs(8165);
    layer1_outputs(6068) <= not(layer0_outputs(935));
    layer1_outputs(6069) <= not(layer0_outputs(3047));
    layer1_outputs(6070) <= not(layer0_outputs(5409));
    layer1_outputs(6071) <= not(layer0_outputs(8538)) or (layer0_outputs(8741));
    layer1_outputs(6072) <= not((layer0_outputs(4428)) and (layer0_outputs(9895)));
    layer1_outputs(6073) <= not((layer0_outputs(752)) and (layer0_outputs(9856)));
    layer1_outputs(6074) <= not(layer0_outputs(6203)) or (layer0_outputs(5774));
    layer1_outputs(6075) <= layer0_outputs(7795);
    layer1_outputs(6076) <= not(layer0_outputs(4454));
    layer1_outputs(6077) <= not(layer0_outputs(4038));
    layer1_outputs(6078) <= not((layer0_outputs(10015)) or (layer0_outputs(9922)));
    layer1_outputs(6079) <= (layer0_outputs(8981)) and not (layer0_outputs(4922));
    layer1_outputs(6080) <= not(layer0_outputs(5659));
    layer1_outputs(6081) <= '1';
    layer1_outputs(6082) <= layer0_outputs(7448);
    layer1_outputs(6083) <= not(layer0_outputs(5772));
    layer1_outputs(6084) <= layer0_outputs(5938);
    layer1_outputs(6085) <= not(layer0_outputs(5182));
    layer1_outputs(6086) <= not(layer0_outputs(8906));
    layer1_outputs(6087) <= not((layer0_outputs(2990)) xor (layer0_outputs(7358)));
    layer1_outputs(6088) <= layer0_outputs(9219);
    layer1_outputs(6089) <= layer0_outputs(4393);
    layer1_outputs(6090) <= layer0_outputs(9900);
    layer1_outputs(6091) <= '1';
    layer1_outputs(6092) <= layer0_outputs(2282);
    layer1_outputs(6093) <= not(layer0_outputs(8492)) or (layer0_outputs(7073));
    layer1_outputs(6094) <= layer0_outputs(1290);
    layer1_outputs(6095) <= (layer0_outputs(8097)) and (layer0_outputs(8094));
    layer1_outputs(6096) <= '1';
    layer1_outputs(6097) <= layer0_outputs(8672);
    layer1_outputs(6098) <= layer0_outputs(1136);
    layer1_outputs(6099) <= (layer0_outputs(9132)) and (layer0_outputs(7517));
    layer1_outputs(6100) <= not(layer0_outputs(5298)) or (layer0_outputs(8385));
    layer1_outputs(6101) <= layer0_outputs(7652);
    layer1_outputs(6102) <= not(layer0_outputs(10160));
    layer1_outputs(6103) <= not(layer0_outputs(2362));
    layer1_outputs(6104) <= not((layer0_outputs(9599)) and (layer0_outputs(1906)));
    layer1_outputs(6105) <= (layer0_outputs(1671)) xor (layer0_outputs(4441));
    layer1_outputs(6106) <= not(layer0_outputs(5077));
    layer1_outputs(6107) <= not(layer0_outputs(5231)) or (layer0_outputs(8523));
    layer1_outputs(6108) <= not(layer0_outputs(9048)) or (layer0_outputs(9538));
    layer1_outputs(6109) <= layer0_outputs(7957);
    layer1_outputs(6110) <= not(layer0_outputs(8138));
    layer1_outputs(6111) <= not(layer0_outputs(6262));
    layer1_outputs(6112) <= layer0_outputs(258);
    layer1_outputs(6113) <= not((layer0_outputs(5963)) and (layer0_outputs(1697)));
    layer1_outputs(6114) <= not(layer0_outputs(4148)) or (layer0_outputs(3976));
    layer1_outputs(6115) <= (layer0_outputs(3651)) or (layer0_outputs(9615));
    layer1_outputs(6116) <= (layer0_outputs(9172)) xor (layer0_outputs(6182));
    layer1_outputs(6117) <= (layer0_outputs(9489)) xor (layer0_outputs(10150));
    layer1_outputs(6118) <= not((layer0_outputs(2722)) or (layer0_outputs(6616)));
    layer1_outputs(6119) <= layer0_outputs(6610);
    layer1_outputs(6120) <= not(layer0_outputs(4507));
    layer1_outputs(6121) <= (layer0_outputs(8334)) and not (layer0_outputs(9668));
    layer1_outputs(6122) <= (layer0_outputs(5420)) and not (layer0_outputs(1679));
    layer1_outputs(6123) <= not((layer0_outputs(2440)) and (layer0_outputs(7277)));
    layer1_outputs(6124) <= (layer0_outputs(6718)) and not (layer0_outputs(1821));
    layer1_outputs(6125) <= (layer0_outputs(4457)) or (layer0_outputs(2184));
    layer1_outputs(6126) <= not(layer0_outputs(7032));
    layer1_outputs(6127) <= '1';
    layer1_outputs(6128) <= (layer0_outputs(5560)) xor (layer0_outputs(3761));
    layer1_outputs(6129) <= (layer0_outputs(5903)) and not (layer0_outputs(1273));
    layer1_outputs(6130) <= not((layer0_outputs(2188)) xor (layer0_outputs(304)));
    layer1_outputs(6131) <= not(layer0_outputs(5119));
    layer1_outputs(6132) <= not(layer0_outputs(3826));
    layer1_outputs(6133) <= not(layer0_outputs(3743));
    layer1_outputs(6134) <= layer0_outputs(7719);
    layer1_outputs(6135) <= (layer0_outputs(7310)) xor (layer0_outputs(2333));
    layer1_outputs(6136) <= not(layer0_outputs(1312));
    layer1_outputs(6137) <= layer0_outputs(5273);
    layer1_outputs(6138) <= (layer0_outputs(8274)) and not (layer0_outputs(426));
    layer1_outputs(6139) <= layer0_outputs(8161);
    layer1_outputs(6140) <= not(layer0_outputs(8068)) or (layer0_outputs(2080));
    layer1_outputs(6141) <= layer0_outputs(1733);
    layer1_outputs(6142) <= '0';
    layer1_outputs(6143) <= (layer0_outputs(6317)) and not (layer0_outputs(762));
    layer1_outputs(6144) <= layer0_outputs(4742);
    layer1_outputs(6145) <= (layer0_outputs(9641)) and not (layer0_outputs(6369));
    layer1_outputs(6146) <= layer0_outputs(4144);
    layer1_outputs(6147) <= not((layer0_outputs(7810)) and (layer0_outputs(5066)));
    layer1_outputs(6148) <= layer0_outputs(6465);
    layer1_outputs(6149) <= not((layer0_outputs(4644)) xor (layer0_outputs(1199)));
    layer1_outputs(6150) <= not(layer0_outputs(3088)) or (layer0_outputs(9183));
    layer1_outputs(6151) <= layer0_outputs(4932);
    layer1_outputs(6152) <= '0';
    layer1_outputs(6153) <= not((layer0_outputs(6945)) and (layer0_outputs(6168)));
    layer1_outputs(6154) <= (layer0_outputs(8354)) or (layer0_outputs(1198));
    layer1_outputs(6155) <= not((layer0_outputs(7099)) or (layer0_outputs(8612)));
    layer1_outputs(6156) <= (layer0_outputs(6684)) or (layer0_outputs(3813));
    layer1_outputs(6157) <= (layer0_outputs(809)) xor (layer0_outputs(9986));
    layer1_outputs(6158) <= layer0_outputs(3241);
    layer1_outputs(6159) <= not(layer0_outputs(3751)) or (layer0_outputs(5751));
    layer1_outputs(6160) <= (layer0_outputs(2775)) and not (layer0_outputs(8233));
    layer1_outputs(6161) <= not(layer0_outputs(9467));
    layer1_outputs(6162) <= not((layer0_outputs(285)) xor (layer0_outputs(1576)));
    layer1_outputs(6163) <= not(layer0_outputs(7700)) or (layer0_outputs(773));
    layer1_outputs(6164) <= not((layer0_outputs(6370)) and (layer0_outputs(6478)));
    layer1_outputs(6165) <= not(layer0_outputs(3542));
    layer1_outputs(6166) <= not((layer0_outputs(2505)) or (layer0_outputs(431)));
    layer1_outputs(6167) <= not((layer0_outputs(7229)) and (layer0_outputs(5291)));
    layer1_outputs(6168) <= not((layer0_outputs(3710)) or (layer0_outputs(4512)));
    layer1_outputs(6169) <= (layer0_outputs(530)) or (layer0_outputs(8331));
    layer1_outputs(6170) <= not((layer0_outputs(3102)) xor (layer0_outputs(2607)));
    layer1_outputs(6171) <= (layer0_outputs(9953)) and not (layer0_outputs(6485));
    layer1_outputs(6172) <= not(layer0_outputs(2660));
    layer1_outputs(6173) <= (layer0_outputs(322)) and (layer0_outputs(2659));
    layer1_outputs(6174) <= layer0_outputs(5230);
    layer1_outputs(6175) <= not(layer0_outputs(1219));
    layer1_outputs(6176) <= not(layer0_outputs(9378)) or (layer0_outputs(4225));
    layer1_outputs(6177) <= not((layer0_outputs(9754)) and (layer0_outputs(4983)));
    layer1_outputs(6178) <= not((layer0_outputs(5199)) or (layer0_outputs(1080)));
    layer1_outputs(6179) <= (layer0_outputs(3700)) and not (layer0_outputs(2642));
    layer1_outputs(6180) <= not(layer0_outputs(6140));
    layer1_outputs(6181) <= not(layer0_outputs(6965)) or (layer0_outputs(10095));
    layer1_outputs(6182) <= not((layer0_outputs(5401)) xor (layer0_outputs(2980)));
    layer1_outputs(6183) <= (layer0_outputs(9572)) and not (layer0_outputs(7535));
    layer1_outputs(6184) <= not(layer0_outputs(8197));
    layer1_outputs(6185) <= (layer0_outputs(7953)) or (layer0_outputs(3923));
    layer1_outputs(6186) <= not(layer0_outputs(5212));
    layer1_outputs(6187) <= (layer0_outputs(674)) and (layer0_outputs(7254));
    layer1_outputs(6188) <= (layer0_outputs(4535)) and not (layer0_outputs(9667));
    layer1_outputs(6189) <= (layer0_outputs(6681)) xor (layer0_outputs(9393));
    layer1_outputs(6190) <= not((layer0_outputs(1767)) and (layer0_outputs(6057)));
    layer1_outputs(6191) <= not((layer0_outputs(5820)) or (layer0_outputs(2889)));
    layer1_outputs(6192) <= not((layer0_outputs(7021)) xor (layer0_outputs(4605)));
    layer1_outputs(6193) <= layer0_outputs(10121);
    layer1_outputs(6194) <= not(layer0_outputs(9832));
    layer1_outputs(6195) <= (layer0_outputs(9776)) or (layer0_outputs(9870));
    layer1_outputs(6196) <= layer0_outputs(7449);
    layer1_outputs(6197) <= not(layer0_outputs(4875));
    layer1_outputs(6198) <= (layer0_outputs(2845)) xor (layer0_outputs(4310));
    layer1_outputs(6199) <= (layer0_outputs(8230)) and not (layer0_outputs(1950));
    layer1_outputs(6200) <= layer0_outputs(6178);
    layer1_outputs(6201) <= (layer0_outputs(4124)) and not (layer0_outputs(8044));
    layer1_outputs(6202) <= layer0_outputs(6000);
    layer1_outputs(6203) <= not((layer0_outputs(2325)) and (layer0_outputs(1508)));
    layer1_outputs(6204) <= (layer0_outputs(6441)) and (layer0_outputs(6848));
    layer1_outputs(6205) <= not(layer0_outputs(1838));
    layer1_outputs(6206) <= not(layer0_outputs(3770));
    layer1_outputs(6207) <= (layer0_outputs(3419)) or (layer0_outputs(6841));
    layer1_outputs(6208) <= '1';
    layer1_outputs(6209) <= not(layer0_outputs(3037));
    layer1_outputs(6210) <= not(layer0_outputs(9983)) or (layer0_outputs(434));
    layer1_outputs(6211) <= layer0_outputs(31);
    layer1_outputs(6212) <= not((layer0_outputs(8746)) and (layer0_outputs(4354)));
    layer1_outputs(6213) <= (layer0_outputs(2005)) and not (layer0_outputs(2320));
    layer1_outputs(6214) <= (layer0_outputs(4236)) or (layer0_outputs(5720));
    layer1_outputs(6215) <= not(layer0_outputs(3037)) or (layer0_outputs(1805));
    layer1_outputs(6216) <= not(layer0_outputs(3588));
    layer1_outputs(6217) <= (layer0_outputs(5440)) xor (layer0_outputs(1880));
    layer1_outputs(6218) <= not((layer0_outputs(9352)) or (layer0_outputs(9735)));
    layer1_outputs(6219) <= layer0_outputs(4930);
    layer1_outputs(6220) <= (layer0_outputs(5471)) and not (layer0_outputs(753));
    layer1_outputs(6221) <= (layer0_outputs(5643)) and not (layer0_outputs(7705));
    layer1_outputs(6222) <= (layer0_outputs(6349)) xor (layer0_outputs(3651));
    layer1_outputs(6223) <= layer0_outputs(4030);
    layer1_outputs(6224) <= '1';
    layer1_outputs(6225) <= not(layer0_outputs(8227));
    layer1_outputs(6226) <= layer0_outputs(5496);
    layer1_outputs(6227) <= '1';
    layer1_outputs(6228) <= layer0_outputs(4712);
    layer1_outputs(6229) <= not(layer0_outputs(7680));
    layer1_outputs(6230) <= not(layer0_outputs(1739));
    layer1_outputs(6231) <= not((layer0_outputs(8921)) xor (layer0_outputs(3939)));
    layer1_outputs(6232) <= not(layer0_outputs(3350));
    layer1_outputs(6233) <= layer0_outputs(8710);
    layer1_outputs(6234) <= not(layer0_outputs(7044)) or (layer0_outputs(1006));
    layer1_outputs(6235) <= not((layer0_outputs(4355)) and (layer0_outputs(1687)));
    layer1_outputs(6236) <= not(layer0_outputs(5828)) or (layer0_outputs(2325));
    layer1_outputs(6237) <= not(layer0_outputs(7461)) or (layer0_outputs(3203));
    layer1_outputs(6238) <= not(layer0_outputs(179));
    layer1_outputs(6239) <= not((layer0_outputs(6522)) and (layer0_outputs(4456)));
    layer1_outputs(6240) <= not(layer0_outputs(4294)) or (layer0_outputs(2705));
    layer1_outputs(6241) <= (layer0_outputs(1954)) and (layer0_outputs(6873));
    layer1_outputs(6242) <= (layer0_outputs(9635)) and not (layer0_outputs(7369));
    layer1_outputs(6243) <= layer0_outputs(3161);
    layer1_outputs(6244) <= not(layer0_outputs(855));
    layer1_outputs(6245) <= not((layer0_outputs(5832)) and (layer0_outputs(9165)));
    layer1_outputs(6246) <= not((layer0_outputs(5200)) or (layer0_outputs(9232)));
    layer1_outputs(6247) <= not(layer0_outputs(7174));
    layer1_outputs(6248) <= (layer0_outputs(3012)) or (layer0_outputs(7005));
    layer1_outputs(6249) <= (layer0_outputs(6866)) or (layer0_outputs(5473));
    layer1_outputs(6250) <= not((layer0_outputs(7975)) xor (layer0_outputs(9959)));
    layer1_outputs(6251) <= (layer0_outputs(5157)) and not (layer0_outputs(5971));
    layer1_outputs(6252) <= (layer0_outputs(6609)) or (layer0_outputs(1962));
    layer1_outputs(6253) <= layer0_outputs(7041);
    layer1_outputs(6254) <= layer0_outputs(5512);
    layer1_outputs(6255) <= not(layer0_outputs(6167));
    layer1_outputs(6256) <= not(layer0_outputs(3959));
    layer1_outputs(6257) <= (layer0_outputs(8909)) xor (layer0_outputs(870));
    layer1_outputs(6258) <= not((layer0_outputs(3145)) xor (layer0_outputs(5057)));
    layer1_outputs(6259) <= not(layer0_outputs(7827)) or (layer0_outputs(1081));
    layer1_outputs(6260) <= not(layer0_outputs(821));
    layer1_outputs(6261) <= not(layer0_outputs(4303));
    layer1_outputs(6262) <= (layer0_outputs(4225)) and (layer0_outputs(4140));
    layer1_outputs(6263) <= layer0_outputs(3451);
    layer1_outputs(6264) <= layer0_outputs(4267);
    layer1_outputs(6265) <= not(layer0_outputs(6491)) or (layer0_outputs(1920));
    layer1_outputs(6266) <= '1';
    layer1_outputs(6267) <= (layer0_outputs(6580)) and (layer0_outputs(7439));
    layer1_outputs(6268) <= layer0_outputs(2874);
    layer1_outputs(6269) <= not(layer0_outputs(229));
    layer1_outputs(6270) <= (layer0_outputs(9621)) xor (layer0_outputs(907));
    layer1_outputs(6271) <= (layer0_outputs(497)) and (layer0_outputs(3565));
    layer1_outputs(6272) <= (layer0_outputs(7384)) and (layer0_outputs(7745));
    layer1_outputs(6273) <= not((layer0_outputs(6181)) xor (layer0_outputs(3842)));
    layer1_outputs(6274) <= (layer0_outputs(769)) or (layer0_outputs(7863));
    layer1_outputs(6275) <= layer0_outputs(2861);
    layer1_outputs(6276) <= not(layer0_outputs(6124)) or (layer0_outputs(1061));
    layer1_outputs(6277) <= not((layer0_outputs(8130)) or (layer0_outputs(8919)));
    layer1_outputs(6278) <= layer0_outputs(8142);
    layer1_outputs(6279) <= layer0_outputs(3380);
    layer1_outputs(6280) <= (layer0_outputs(3948)) xor (layer0_outputs(6734));
    layer1_outputs(6281) <= not(layer0_outputs(3398));
    layer1_outputs(6282) <= layer0_outputs(7386);
    layer1_outputs(6283) <= not(layer0_outputs(131));
    layer1_outputs(6284) <= not(layer0_outputs(7285));
    layer1_outputs(6285) <= not((layer0_outputs(9678)) or (layer0_outputs(10124)));
    layer1_outputs(6286) <= not(layer0_outputs(3862));
    layer1_outputs(6287) <= (layer0_outputs(7221)) and not (layer0_outputs(2403));
    layer1_outputs(6288) <= layer0_outputs(6434);
    layer1_outputs(6289) <= layer0_outputs(3145);
    layer1_outputs(6290) <= not(layer0_outputs(3630));
    layer1_outputs(6291) <= '1';
    layer1_outputs(6292) <= not((layer0_outputs(2032)) and (layer0_outputs(3445)));
    layer1_outputs(6293) <= not((layer0_outputs(2186)) or (layer0_outputs(5704)));
    layer1_outputs(6294) <= not(layer0_outputs(5188));
    layer1_outputs(6295) <= not(layer0_outputs(408)) or (layer0_outputs(1020));
    layer1_outputs(6296) <= not(layer0_outputs(974));
    layer1_outputs(6297) <= not(layer0_outputs(10127)) or (layer0_outputs(4545));
    layer1_outputs(6298) <= (layer0_outputs(199)) or (layer0_outputs(7462));
    layer1_outputs(6299) <= (layer0_outputs(2787)) or (layer0_outputs(6375));
    layer1_outputs(6300) <= not(layer0_outputs(4412)) or (layer0_outputs(503));
    layer1_outputs(6301) <= (layer0_outputs(5095)) and (layer0_outputs(8408));
    layer1_outputs(6302) <= not(layer0_outputs(7972)) or (layer0_outputs(1294));
    layer1_outputs(6303) <= not(layer0_outputs(7753));
    layer1_outputs(6304) <= not(layer0_outputs(8485));
    layer1_outputs(6305) <= layer0_outputs(9322);
    layer1_outputs(6306) <= not(layer0_outputs(3559)) or (layer0_outputs(3166));
    layer1_outputs(6307) <= not(layer0_outputs(9000));
    layer1_outputs(6308) <= not(layer0_outputs(7595)) or (layer0_outputs(2183));
    layer1_outputs(6309) <= layer0_outputs(4026);
    layer1_outputs(6310) <= (layer0_outputs(6224)) or (layer0_outputs(1907));
    layer1_outputs(6311) <= (layer0_outputs(4523)) xor (layer0_outputs(908));
    layer1_outputs(6312) <= (layer0_outputs(4734)) or (layer0_outputs(3856));
    layer1_outputs(6313) <= layer0_outputs(3507);
    layer1_outputs(6314) <= (layer0_outputs(7451)) or (layer0_outputs(5820));
    layer1_outputs(6315) <= layer0_outputs(8504);
    layer1_outputs(6316) <= layer0_outputs(4610);
    layer1_outputs(6317) <= not(layer0_outputs(9340));
    layer1_outputs(6318) <= layer0_outputs(7829);
    layer1_outputs(6319) <= not((layer0_outputs(6147)) and (layer0_outputs(4409)));
    layer1_outputs(6320) <= layer0_outputs(7617);
    layer1_outputs(6321) <= not(layer0_outputs(6259));
    layer1_outputs(6322) <= layer0_outputs(9115);
    layer1_outputs(6323) <= layer0_outputs(10118);
    layer1_outputs(6324) <= not(layer0_outputs(1379));
    layer1_outputs(6325) <= not(layer0_outputs(3685)) or (layer0_outputs(3047));
    layer1_outputs(6326) <= not(layer0_outputs(2766));
    layer1_outputs(6327) <= layer0_outputs(6952);
    layer1_outputs(6328) <= not((layer0_outputs(5208)) or (layer0_outputs(4432)));
    layer1_outputs(6329) <= not((layer0_outputs(3457)) xor (layer0_outputs(2753)));
    layer1_outputs(6330) <= not(layer0_outputs(10165)) or (layer0_outputs(1943));
    layer1_outputs(6331) <= not(layer0_outputs(1347)) or (layer0_outputs(7351));
    layer1_outputs(6332) <= (layer0_outputs(2514)) and not (layer0_outputs(5070));
    layer1_outputs(6333) <= (layer0_outputs(7054)) and not (layer0_outputs(2348));
    layer1_outputs(6334) <= not(layer0_outputs(927));
    layer1_outputs(6335) <= not((layer0_outputs(2663)) and (layer0_outputs(5544)));
    layer1_outputs(6336) <= not((layer0_outputs(1107)) or (layer0_outputs(3342)));
    layer1_outputs(6337) <= not((layer0_outputs(3718)) and (layer0_outputs(1183)));
    layer1_outputs(6338) <= (layer0_outputs(1174)) and not (layer0_outputs(8727));
    layer1_outputs(6339) <= not(layer0_outputs(4725));
    layer1_outputs(6340) <= not(layer0_outputs(5591));
    layer1_outputs(6341) <= not(layer0_outputs(402)) or (layer0_outputs(5394));
    layer1_outputs(6342) <= not((layer0_outputs(2587)) xor (layer0_outputs(8141)));
    layer1_outputs(6343) <= layer0_outputs(2183);
    layer1_outputs(6344) <= not(layer0_outputs(8873));
    layer1_outputs(6345) <= not(layer0_outputs(2265));
    layer1_outputs(6346) <= (layer0_outputs(9527)) and not (layer0_outputs(2496));
    layer1_outputs(6347) <= not(layer0_outputs(516)) or (layer0_outputs(8509));
    layer1_outputs(6348) <= not(layer0_outputs(2308));
    layer1_outputs(6349) <= not(layer0_outputs(2268));
    layer1_outputs(6350) <= not(layer0_outputs(4981));
    layer1_outputs(6351) <= not((layer0_outputs(9852)) or (layer0_outputs(7958)));
    layer1_outputs(6352) <= (layer0_outputs(5805)) and not (layer0_outputs(5196));
    layer1_outputs(6353) <= not(layer0_outputs(4244));
    layer1_outputs(6354) <= not(layer0_outputs(5984)) or (layer0_outputs(8875));
    layer1_outputs(6355) <= not(layer0_outputs(6942));
    layer1_outputs(6356) <= (layer0_outputs(6860)) and (layer0_outputs(9223));
    layer1_outputs(6357) <= not(layer0_outputs(5993));
    layer1_outputs(6358) <= (layer0_outputs(10112)) or (layer0_outputs(777));
    layer1_outputs(6359) <= (layer0_outputs(1612)) and not (layer0_outputs(4235));
    layer1_outputs(6360) <= (layer0_outputs(4126)) and not (layer0_outputs(116));
    layer1_outputs(6361) <= (layer0_outputs(5816)) and not (layer0_outputs(4999));
    layer1_outputs(6362) <= (layer0_outputs(896)) xor (layer0_outputs(3861));
    layer1_outputs(6363) <= not((layer0_outputs(6330)) and (layer0_outputs(7738)));
    layer1_outputs(6364) <= not((layer0_outputs(4518)) and (layer0_outputs(82)));
    layer1_outputs(6365) <= not(layer0_outputs(3609)) or (layer0_outputs(6197));
    layer1_outputs(6366) <= not((layer0_outputs(9742)) xor (layer0_outputs(4841)));
    layer1_outputs(6367) <= not(layer0_outputs(6111)) or (layer0_outputs(2948));
    layer1_outputs(6368) <= not(layer0_outputs(4680));
    layer1_outputs(6369) <= not(layer0_outputs(7962));
    layer1_outputs(6370) <= not(layer0_outputs(9021)) or (layer0_outputs(6899));
    layer1_outputs(6371) <= (layer0_outputs(1930)) and not (layer0_outputs(8885));
    layer1_outputs(6372) <= (layer0_outputs(9477)) and not (layer0_outputs(9146));
    layer1_outputs(6373) <= not(layer0_outputs(4971));
    layer1_outputs(6374) <= not((layer0_outputs(1527)) or (layer0_outputs(4456)));
    layer1_outputs(6375) <= not(layer0_outputs(9359)) or (layer0_outputs(120));
    layer1_outputs(6376) <= not(layer0_outputs(2302)) or (layer0_outputs(2779));
    layer1_outputs(6377) <= (layer0_outputs(7331)) and not (layer0_outputs(3669));
    layer1_outputs(6378) <= (layer0_outputs(5386)) or (layer0_outputs(6947));
    layer1_outputs(6379) <= (layer0_outputs(2859)) and (layer0_outputs(348));
    layer1_outputs(6380) <= (layer0_outputs(3295)) and (layer0_outputs(9244));
    layer1_outputs(6381) <= not((layer0_outputs(10060)) xor (layer0_outputs(48)));
    layer1_outputs(6382) <= not(layer0_outputs(2549)) or (layer0_outputs(6861));
    layer1_outputs(6383) <= (layer0_outputs(513)) xor (layer0_outputs(3531));
    layer1_outputs(6384) <= layer0_outputs(7056);
    layer1_outputs(6385) <= (layer0_outputs(9444)) and not (layer0_outputs(327));
    layer1_outputs(6386) <= not(layer0_outputs(8928));
    layer1_outputs(6387) <= layer0_outputs(7592);
    layer1_outputs(6388) <= not((layer0_outputs(9255)) and (layer0_outputs(4588)));
    layer1_outputs(6389) <= not(layer0_outputs(9238));
    layer1_outputs(6390) <= not(layer0_outputs(1783));
    layer1_outputs(6391) <= layer0_outputs(907);
    layer1_outputs(6392) <= '1';
    layer1_outputs(6393) <= '0';
    layer1_outputs(6394) <= not(layer0_outputs(5295));
    layer1_outputs(6395) <= (layer0_outputs(4137)) and not (layer0_outputs(1043));
    layer1_outputs(6396) <= (layer0_outputs(5058)) or (layer0_outputs(3623));
    layer1_outputs(6397) <= not((layer0_outputs(4322)) and (layer0_outputs(8999)));
    layer1_outputs(6398) <= not(layer0_outputs(460)) or (layer0_outputs(1417));
    layer1_outputs(6399) <= (layer0_outputs(2047)) and not (layer0_outputs(649));
    layer1_outputs(6400) <= (layer0_outputs(815)) and (layer0_outputs(46));
    layer1_outputs(6401) <= layer0_outputs(598);
    layer1_outputs(6402) <= layer0_outputs(1311);
    layer1_outputs(6403) <= not((layer0_outputs(9001)) xor (layer0_outputs(1164)));
    layer1_outputs(6404) <= (layer0_outputs(6417)) and not (layer0_outputs(2133));
    layer1_outputs(6405) <= not(layer0_outputs(5045)) or (layer0_outputs(2420));
    layer1_outputs(6406) <= not(layer0_outputs(7157));
    layer1_outputs(6407) <= not(layer0_outputs(8576));
    layer1_outputs(6408) <= not(layer0_outputs(8896)) or (layer0_outputs(10037));
    layer1_outputs(6409) <= (layer0_outputs(6788)) or (layer0_outputs(1204));
    layer1_outputs(6410) <= (layer0_outputs(7392)) or (layer0_outputs(4767));
    layer1_outputs(6411) <= not(layer0_outputs(4408)) or (layer0_outputs(9136));
    layer1_outputs(6412) <= not((layer0_outputs(3412)) or (layer0_outputs(1197)));
    layer1_outputs(6413) <= layer0_outputs(2745);
    layer1_outputs(6414) <= layer0_outputs(596);
    layer1_outputs(6415) <= layer0_outputs(1106);
    layer1_outputs(6416) <= layer0_outputs(9891);
    layer1_outputs(6417) <= '0';
    layer1_outputs(6418) <= layer0_outputs(8536);
    layer1_outputs(6419) <= layer0_outputs(3000);
    layer1_outputs(6420) <= not((layer0_outputs(5749)) or (layer0_outputs(8832)));
    layer1_outputs(6421) <= not(layer0_outputs(2695));
    layer1_outputs(6422) <= not(layer0_outputs(1665));
    layer1_outputs(6423) <= not(layer0_outputs(9228)) or (layer0_outputs(1140));
    layer1_outputs(6424) <= not(layer0_outputs(3838));
    layer1_outputs(6425) <= not(layer0_outputs(8749));
    layer1_outputs(6426) <= not(layer0_outputs(4909));
    layer1_outputs(6427) <= layer0_outputs(5017);
    layer1_outputs(6428) <= not((layer0_outputs(5389)) or (layer0_outputs(10075)));
    layer1_outputs(6429) <= layer0_outputs(8004);
    layer1_outputs(6430) <= layer0_outputs(1553);
    layer1_outputs(6431) <= not((layer0_outputs(8661)) and (layer0_outputs(2674)));
    layer1_outputs(6432) <= layer0_outputs(6454);
    layer1_outputs(6433) <= not((layer0_outputs(6294)) xor (layer0_outputs(5964)));
    layer1_outputs(6434) <= not(layer0_outputs(795));
    layer1_outputs(6435) <= not(layer0_outputs(9848));
    layer1_outputs(6436) <= layer0_outputs(7096);
    layer1_outputs(6437) <= layer0_outputs(7440);
    layer1_outputs(6438) <= not(layer0_outputs(3125)) or (layer0_outputs(1708));
    layer1_outputs(6439) <= not(layer0_outputs(1660)) or (layer0_outputs(797));
    layer1_outputs(6440) <= not((layer0_outputs(1596)) xor (layer0_outputs(8722)));
    layer1_outputs(6441) <= not(layer0_outputs(4012)) or (layer0_outputs(6051));
    layer1_outputs(6442) <= '1';
    layer1_outputs(6443) <= not((layer0_outputs(719)) and (layer0_outputs(1713)));
    layer1_outputs(6444) <= not((layer0_outputs(3186)) and (layer0_outputs(8394)));
    layer1_outputs(6445) <= not((layer0_outputs(9175)) or (layer0_outputs(447)));
    layer1_outputs(6446) <= not((layer0_outputs(2982)) xor (layer0_outputs(4420)));
    layer1_outputs(6447) <= not((layer0_outputs(4129)) and (layer0_outputs(9684)));
    layer1_outputs(6448) <= layer0_outputs(9441);
    layer1_outputs(6449) <= (layer0_outputs(8052)) or (layer0_outputs(7045));
    layer1_outputs(6450) <= layer0_outputs(553);
    layer1_outputs(6451) <= layer0_outputs(3410);
    layer1_outputs(6452) <= not((layer0_outputs(9976)) or (layer0_outputs(297)));
    layer1_outputs(6453) <= layer0_outputs(7105);
    layer1_outputs(6454) <= not(layer0_outputs(7919)) or (layer0_outputs(9362));
    layer1_outputs(6455) <= (layer0_outputs(6832)) and not (layer0_outputs(5783));
    layer1_outputs(6456) <= (layer0_outputs(1594)) and (layer0_outputs(5416));
    layer1_outputs(6457) <= (layer0_outputs(3127)) and (layer0_outputs(5097));
    layer1_outputs(6458) <= not(layer0_outputs(9482)) or (layer0_outputs(852));
    layer1_outputs(6459) <= not(layer0_outputs(1029));
    layer1_outputs(6460) <= not(layer0_outputs(7554)) or (layer0_outputs(498));
    layer1_outputs(6461) <= (layer0_outputs(6743)) and (layer0_outputs(1806));
    layer1_outputs(6462) <= not(layer0_outputs(3292));
    layer1_outputs(6463) <= not(layer0_outputs(9186));
    layer1_outputs(6464) <= (layer0_outputs(2235)) and not (layer0_outputs(2431));
    layer1_outputs(6465) <= (layer0_outputs(6808)) and not (layer0_outputs(3604));
    layer1_outputs(6466) <= (layer0_outputs(9413)) and not (layer0_outputs(5518));
    layer1_outputs(6467) <= layer0_outputs(7388);
    layer1_outputs(6468) <= layer0_outputs(7185);
    layer1_outputs(6469) <= layer0_outputs(1850);
    layer1_outputs(6470) <= layer0_outputs(1906);
    layer1_outputs(6471) <= (layer0_outputs(8093)) or (layer0_outputs(5858));
    layer1_outputs(6472) <= '0';
    layer1_outputs(6473) <= not(layer0_outputs(2132));
    layer1_outputs(6474) <= (layer0_outputs(6473)) or (layer0_outputs(6636));
    layer1_outputs(6475) <= (layer0_outputs(3520)) and (layer0_outputs(6991));
    layer1_outputs(6476) <= not(layer0_outputs(6613)) or (layer0_outputs(3612));
    layer1_outputs(6477) <= not(layer0_outputs(177)) or (layer0_outputs(2374));
    layer1_outputs(6478) <= layer0_outputs(1476);
    layer1_outputs(6479) <= layer0_outputs(7704);
    layer1_outputs(6480) <= not(layer0_outputs(8952)) or (layer0_outputs(2405));
    layer1_outputs(6481) <= layer0_outputs(8595);
    layer1_outputs(6482) <= not(layer0_outputs(7230)) or (layer0_outputs(4496));
    layer1_outputs(6483) <= (layer0_outputs(7899)) or (layer0_outputs(496));
    layer1_outputs(6484) <= layer0_outputs(4163);
    layer1_outputs(6485) <= layer0_outputs(857);
    layer1_outputs(6486) <= not(layer0_outputs(1514));
    layer1_outputs(6487) <= not(layer0_outputs(4785));
    layer1_outputs(6488) <= layer0_outputs(10205);
    layer1_outputs(6489) <= not(layer0_outputs(1815));
    layer1_outputs(6490) <= not((layer0_outputs(7104)) or (layer0_outputs(3117)));
    layer1_outputs(6491) <= layer0_outputs(4022);
    layer1_outputs(6492) <= not(layer0_outputs(1380)) or (layer0_outputs(9277));
    layer1_outputs(6493) <= not((layer0_outputs(9183)) or (layer0_outputs(2606)));
    layer1_outputs(6494) <= (layer0_outputs(3602)) and not (layer0_outputs(4452));
    layer1_outputs(6495) <= layer0_outputs(10193);
    layer1_outputs(6496) <= not((layer0_outputs(3192)) and (layer0_outputs(4631)));
    layer1_outputs(6497) <= (layer0_outputs(647)) or (layer0_outputs(8070));
    layer1_outputs(6498) <= layer0_outputs(6363);
    layer1_outputs(6499) <= layer0_outputs(6540);
    layer1_outputs(6500) <= not(layer0_outputs(2552));
    layer1_outputs(6501) <= layer0_outputs(2713);
    layer1_outputs(6502) <= not((layer0_outputs(3963)) or (layer0_outputs(838)));
    layer1_outputs(6503) <= layer0_outputs(5185);
    layer1_outputs(6504) <= layer0_outputs(3110);
    layer1_outputs(6505) <= (layer0_outputs(7744)) and not (layer0_outputs(1966));
    layer1_outputs(6506) <= not(layer0_outputs(1121));
    layer1_outputs(6507) <= not(layer0_outputs(3144));
    layer1_outputs(6508) <= (layer0_outputs(476)) xor (layer0_outputs(1662));
    layer1_outputs(6509) <= not((layer0_outputs(1871)) xor (layer0_outputs(2593)));
    layer1_outputs(6510) <= not(layer0_outputs(7867));
    layer1_outputs(6511) <= layer0_outputs(3822);
    layer1_outputs(6512) <= layer0_outputs(595);
    layer1_outputs(6513) <= (layer0_outputs(2612)) and not (layer0_outputs(6940));
    layer1_outputs(6514) <= (layer0_outputs(6298)) and not (layer0_outputs(2391));
    layer1_outputs(6515) <= layer0_outputs(9329);
    layer1_outputs(6516) <= not((layer0_outputs(5555)) or (layer0_outputs(7881)));
    layer1_outputs(6517) <= (layer0_outputs(7232)) and not (layer0_outputs(1325));
    layer1_outputs(6518) <= not(layer0_outputs(5213));
    layer1_outputs(6519) <= not(layer0_outputs(2796));
    layer1_outputs(6520) <= layer0_outputs(8664);
    layer1_outputs(6521) <= layer0_outputs(5351);
    layer1_outputs(6522) <= not((layer0_outputs(310)) or (layer0_outputs(8876)));
    layer1_outputs(6523) <= not(layer0_outputs(4331)) or (layer0_outputs(5587));
    layer1_outputs(6524) <= layer0_outputs(8424);
    layer1_outputs(6525) <= (layer0_outputs(373)) and (layer0_outputs(793));
    layer1_outputs(6526) <= not((layer0_outputs(4766)) and (layer0_outputs(1477)));
    layer1_outputs(6527) <= layer0_outputs(4560);
    layer1_outputs(6528) <= (layer0_outputs(585)) and not (layer0_outputs(6824));
    layer1_outputs(6529) <= not(layer0_outputs(3752));
    layer1_outputs(6530) <= not((layer0_outputs(2277)) xor (layer0_outputs(2660)));
    layer1_outputs(6531) <= layer0_outputs(5848);
    layer1_outputs(6532) <= (layer0_outputs(8453)) or (layer0_outputs(1657));
    layer1_outputs(6533) <= not((layer0_outputs(4042)) xor (layer0_outputs(7103)));
    layer1_outputs(6534) <= not(layer0_outputs(5763));
    layer1_outputs(6535) <= not(layer0_outputs(7609)) or (layer0_outputs(7427));
    layer1_outputs(6536) <= (layer0_outputs(9332)) and (layer0_outputs(9114));
    layer1_outputs(6537) <= (layer0_outputs(10188)) and not (layer0_outputs(2565));
    layer1_outputs(6538) <= not(layer0_outputs(227));
    layer1_outputs(6539) <= not(layer0_outputs(925));
    layer1_outputs(6540) <= layer0_outputs(79);
    layer1_outputs(6541) <= layer0_outputs(2457);
    layer1_outputs(6542) <= (layer0_outputs(7175)) and not (layer0_outputs(2562));
    layer1_outputs(6543) <= (layer0_outputs(6993)) and not (layer0_outputs(225));
    layer1_outputs(6544) <= (layer0_outputs(8353)) xor (layer0_outputs(3312));
    layer1_outputs(6545) <= (layer0_outputs(9077)) xor (layer0_outputs(6975));
    layer1_outputs(6546) <= layer0_outputs(4083);
    layer1_outputs(6547) <= layer0_outputs(4025);
    layer1_outputs(6548) <= not((layer0_outputs(5006)) and (layer0_outputs(9548)));
    layer1_outputs(6549) <= layer0_outputs(8780);
    layer1_outputs(6550) <= (layer0_outputs(3388)) and (layer0_outputs(2747));
    layer1_outputs(6551) <= not(layer0_outputs(9065));
    layer1_outputs(6552) <= layer0_outputs(4252);
    layer1_outputs(6553) <= (layer0_outputs(2258)) and (layer0_outputs(9598));
    layer1_outputs(6554) <= (layer0_outputs(5788)) or (layer0_outputs(1229));
    layer1_outputs(6555) <= (layer0_outputs(5655)) and not (layer0_outputs(8575));
    layer1_outputs(6556) <= layer0_outputs(1466);
    layer1_outputs(6557) <= not(layer0_outputs(9869)) or (layer0_outputs(9625));
    layer1_outputs(6558) <= not((layer0_outputs(9388)) xor (layer0_outputs(3233)));
    layer1_outputs(6559) <= (layer0_outputs(4241)) or (layer0_outputs(8886));
    layer1_outputs(6560) <= '0';
    layer1_outputs(6561) <= (layer0_outputs(8506)) or (layer0_outputs(6258));
    layer1_outputs(6562) <= not((layer0_outputs(1413)) and (layer0_outputs(7600)));
    layer1_outputs(6563) <= (layer0_outputs(8501)) or (layer0_outputs(4253));
    layer1_outputs(6564) <= layer0_outputs(7444);
    layer1_outputs(6565) <= '0';
    layer1_outputs(6566) <= (layer0_outputs(7598)) or (layer0_outputs(2617));
    layer1_outputs(6567) <= not(layer0_outputs(254));
    layer1_outputs(6568) <= not((layer0_outputs(6592)) xor (layer0_outputs(6670)));
    layer1_outputs(6569) <= not(layer0_outputs(76));
    layer1_outputs(6570) <= not(layer0_outputs(1800)) or (layer0_outputs(9048));
    layer1_outputs(6571) <= layer0_outputs(638);
    layer1_outputs(6572) <= not((layer0_outputs(2512)) and (layer0_outputs(5505)));
    layer1_outputs(6573) <= (layer0_outputs(4091)) and not (layer0_outputs(7343));
    layer1_outputs(6574) <= not((layer0_outputs(9555)) and (layer0_outputs(4299)));
    layer1_outputs(6575) <= layer0_outputs(8143);
    layer1_outputs(6576) <= (layer0_outputs(9956)) and (layer0_outputs(3314));
    layer1_outputs(6577) <= (layer0_outputs(1802)) or (layer0_outputs(9599));
    layer1_outputs(6578) <= (layer0_outputs(4206)) and not (layer0_outputs(732));
    layer1_outputs(6579) <= not(layer0_outputs(9070));
    layer1_outputs(6580) <= layer0_outputs(10143);
    layer1_outputs(6581) <= (layer0_outputs(8930)) or (layer0_outputs(2246));
    layer1_outputs(6582) <= not(layer0_outputs(6210)) or (layer0_outputs(7309));
    layer1_outputs(6583) <= not((layer0_outputs(3231)) or (layer0_outputs(109)));
    layer1_outputs(6584) <= not(layer0_outputs(4670)) or (layer0_outputs(4639));
    layer1_outputs(6585) <= layer0_outputs(8838);
    layer1_outputs(6586) <= not((layer0_outputs(4894)) and (layer0_outputs(9659)));
    layer1_outputs(6587) <= (layer0_outputs(9963)) xor (layer0_outputs(6126));
    layer1_outputs(6588) <= layer0_outputs(1580);
    layer1_outputs(6589) <= layer0_outputs(7092);
    layer1_outputs(6590) <= not((layer0_outputs(4531)) or (layer0_outputs(253)));
    layer1_outputs(6591) <= layer0_outputs(18);
    layer1_outputs(6592) <= not(layer0_outputs(2395));
    layer1_outputs(6593) <= (layer0_outputs(3644)) and not (layer0_outputs(6050));
    layer1_outputs(6594) <= not((layer0_outputs(2438)) or (layer0_outputs(6103)));
    layer1_outputs(6595) <= layer0_outputs(8543);
    layer1_outputs(6596) <= not(layer0_outputs(8017)) or (layer0_outputs(4077));
    layer1_outputs(6597) <= not(layer0_outputs(1358));
    layer1_outputs(6598) <= (layer0_outputs(7078)) and (layer0_outputs(1395));
    layer1_outputs(6599) <= not((layer0_outputs(3371)) and (layer0_outputs(9493)));
    layer1_outputs(6600) <= not(layer0_outputs(5300));
    layer1_outputs(6601) <= not((layer0_outputs(2825)) or (layer0_outputs(8820)));
    layer1_outputs(6602) <= (layer0_outputs(7239)) or (layer0_outputs(1636));
    layer1_outputs(6603) <= layer0_outputs(8878);
    layer1_outputs(6604) <= not(layer0_outputs(2541));
    layer1_outputs(6605) <= not(layer0_outputs(6459));
    layer1_outputs(6606) <= not(layer0_outputs(7891));
    layer1_outputs(6607) <= (layer0_outputs(6394)) and not (layer0_outputs(3683));
    layer1_outputs(6608) <= (layer0_outputs(3148)) xor (layer0_outputs(9930));
    layer1_outputs(6609) <= (layer0_outputs(2446)) or (layer0_outputs(2007));
    layer1_outputs(6610) <= not(layer0_outputs(4730));
    layer1_outputs(6611) <= not(layer0_outputs(3100));
    layer1_outputs(6612) <= not(layer0_outputs(6830));
    layer1_outputs(6613) <= (layer0_outputs(8233)) or (layer0_outputs(2495));
    layer1_outputs(6614) <= not(layer0_outputs(8753));
    layer1_outputs(6615) <= not((layer0_outputs(5925)) and (layer0_outputs(4016)));
    layer1_outputs(6616) <= layer0_outputs(4157);
    layer1_outputs(6617) <= (layer0_outputs(5902)) xor (layer0_outputs(5837));
    layer1_outputs(6618) <= not(layer0_outputs(3596));
    layer1_outputs(6619) <= layer0_outputs(7032);
    layer1_outputs(6620) <= not((layer0_outputs(119)) xor (layer0_outputs(7009)));
    layer1_outputs(6621) <= layer0_outputs(10118);
    layer1_outputs(6622) <= '0';
    layer1_outputs(6623) <= not((layer0_outputs(5473)) or (layer0_outputs(2707)));
    layer1_outputs(6624) <= not((layer0_outputs(2086)) and (layer0_outputs(9589)));
    layer1_outputs(6625) <= layer0_outputs(6084);
    layer1_outputs(6626) <= not(layer0_outputs(1118)) or (layer0_outputs(4130));
    layer1_outputs(6627) <= layer0_outputs(7172);
    layer1_outputs(6628) <= layer0_outputs(9755);
    layer1_outputs(6629) <= (layer0_outputs(2775)) xor (layer0_outputs(3026));
    layer1_outputs(6630) <= layer0_outputs(2081);
    layer1_outputs(6631) <= not(layer0_outputs(5770)) or (layer0_outputs(5582));
    layer1_outputs(6632) <= not(layer0_outputs(615));
    layer1_outputs(6633) <= not((layer0_outputs(6714)) or (layer0_outputs(7752)));
    layer1_outputs(6634) <= not((layer0_outputs(6806)) xor (layer0_outputs(1241)));
    layer1_outputs(6635) <= (layer0_outputs(2159)) and (layer0_outputs(5588));
    layer1_outputs(6636) <= (layer0_outputs(7002)) and not (layer0_outputs(4806));
    layer1_outputs(6637) <= not((layer0_outputs(9144)) and (layer0_outputs(3548)));
    layer1_outputs(6638) <= not(layer0_outputs(9919));
    layer1_outputs(6639) <= (layer0_outputs(4244)) or (layer0_outputs(9764));
    layer1_outputs(6640) <= layer0_outputs(4367);
    layer1_outputs(6641) <= layer0_outputs(3413);
    layer1_outputs(6642) <= not((layer0_outputs(1322)) and (layer0_outputs(2209)));
    layer1_outputs(6643) <= layer0_outputs(1172);
    layer1_outputs(6644) <= (layer0_outputs(3178)) or (layer0_outputs(3460));
    layer1_outputs(6645) <= (layer0_outputs(4000)) and not (layer0_outputs(3590));
    layer1_outputs(6646) <= not((layer0_outputs(9503)) or (layer0_outputs(9858)));
    layer1_outputs(6647) <= '0';
    layer1_outputs(6648) <= not(layer0_outputs(2304));
    layer1_outputs(6649) <= layer0_outputs(1718);
    layer1_outputs(6650) <= (layer0_outputs(4873)) and (layer0_outputs(2815));
    layer1_outputs(6651) <= layer0_outputs(2419);
    layer1_outputs(6652) <= layer0_outputs(5453);
    layer1_outputs(6653) <= (layer0_outputs(6336)) and (layer0_outputs(8689));
    layer1_outputs(6654) <= not((layer0_outputs(5136)) and (layer0_outputs(8503)));
    layer1_outputs(6655) <= (layer0_outputs(568)) xor (layer0_outputs(3975));
    layer1_outputs(6656) <= layer0_outputs(4281);
    layer1_outputs(6657) <= not((layer0_outputs(2485)) and (layer0_outputs(4320)));
    layer1_outputs(6658) <= not(layer0_outputs(5492));
    layer1_outputs(6659) <= not(layer0_outputs(6257));
    layer1_outputs(6660) <= not((layer0_outputs(7464)) xor (layer0_outputs(4625)));
    layer1_outputs(6661) <= (layer0_outputs(6123)) and (layer0_outputs(6222));
    layer1_outputs(6662) <= '0';
    layer1_outputs(6663) <= not((layer0_outputs(8331)) xor (layer0_outputs(3982)));
    layer1_outputs(6664) <= not(layer0_outputs(6898));
    layer1_outputs(6665) <= (layer0_outputs(7923)) and not (layer0_outputs(8880));
    layer1_outputs(6666) <= layer0_outputs(3740);
    layer1_outputs(6667) <= (layer0_outputs(1989)) and not (layer0_outputs(6523));
    layer1_outputs(6668) <= not(layer0_outputs(4341));
    layer1_outputs(6669) <= (layer0_outputs(7482)) and not (layer0_outputs(378));
    layer1_outputs(6670) <= not(layer0_outputs(1522));
    layer1_outputs(6671) <= layer0_outputs(1425);
    layer1_outputs(6672) <= (layer0_outputs(10187)) and (layer0_outputs(2232));
    layer1_outputs(6673) <= (layer0_outputs(1329)) or (layer0_outputs(9329));
    layer1_outputs(6674) <= (layer0_outputs(5133)) and not (layer0_outputs(3516));
    layer1_outputs(6675) <= (layer0_outputs(8384)) and not (layer0_outputs(2114));
    layer1_outputs(6676) <= (layer0_outputs(6912)) or (layer0_outputs(5503));
    layer1_outputs(6677) <= not(layer0_outputs(5867));
    layer1_outputs(6678) <= (layer0_outputs(10210)) and not (layer0_outputs(5008));
    layer1_outputs(6679) <= (layer0_outputs(229)) xor (layer0_outputs(9540));
    layer1_outputs(6680) <= not(layer0_outputs(2510));
    layer1_outputs(6681) <= not(layer0_outputs(3227)) or (layer0_outputs(3427));
    layer1_outputs(6682) <= not((layer0_outputs(1957)) and (layer0_outputs(2061)));
    layer1_outputs(6683) <= layer0_outputs(5314);
    layer1_outputs(6684) <= (layer0_outputs(2535)) and not (layer0_outputs(8657));
    layer1_outputs(6685) <= (layer0_outputs(6329)) or (layer0_outputs(2052));
    layer1_outputs(6686) <= not(layer0_outputs(391));
    layer1_outputs(6687) <= layer0_outputs(5281);
    layer1_outputs(6688) <= not(layer0_outputs(6496));
    layer1_outputs(6689) <= '1';
    layer1_outputs(6690) <= not(layer0_outputs(7488));
    layer1_outputs(6691) <= not(layer0_outputs(7976));
    layer1_outputs(6692) <= (layer0_outputs(8813)) or (layer0_outputs(189));
    layer1_outputs(6693) <= not((layer0_outputs(2758)) or (layer0_outputs(7199)));
    layer1_outputs(6694) <= not(layer0_outputs(7839));
    layer1_outputs(6695) <= not(layer0_outputs(5302)) or (layer0_outputs(5122));
    layer1_outputs(6696) <= not((layer0_outputs(6515)) xor (layer0_outputs(9923)));
    layer1_outputs(6697) <= (layer0_outputs(380)) and (layer0_outputs(5786));
    layer1_outputs(6698) <= layer0_outputs(286);
    layer1_outputs(6699) <= not((layer0_outputs(6731)) or (layer0_outputs(4230)));
    layer1_outputs(6700) <= '1';
    layer1_outputs(6701) <= layer0_outputs(3953);
    layer1_outputs(6702) <= '0';
    layer1_outputs(6703) <= not(layer0_outputs(5777));
    layer1_outputs(6704) <= (layer0_outputs(5981)) and not (layer0_outputs(1234));
    layer1_outputs(6705) <= not((layer0_outputs(4166)) xor (layer0_outputs(7616)));
    layer1_outputs(6706) <= layer0_outputs(4704);
    layer1_outputs(6707) <= not(layer0_outputs(6348));
    layer1_outputs(6708) <= not((layer0_outputs(2832)) xor (layer0_outputs(4382)));
    layer1_outputs(6709) <= not(layer0_outputs(9653)) or (layer0_outputs(10081));
    layer1_outputs(6710) <= layer0_outputs(3901);
    layer1_outputs(6711) <= layer0_outputs(8540);
    layer1_outputs(6712) <= not(layer0_outputs(922)) or (layer0_outputs(5916));
    layer1_outputs(6713) <= (layer0_outputs(1308)) xor (layer0_outputs(4103));
    layer1_outputs(6714) <= '1';
    layer1_outputs(6715) <= not(layer0_outputs(9884));
    layer1_outputs(6716) <= (layer0_outputs(3144)) xor (layer0_outputs(2633));
    layer1_outputs(6717) <= (layer0_outputs(9748)) and (layer0_outputs(2979));
    layer1_outputs(6718) <= not(layer0_outputs(7431)) or (layer0_outputs(1400));
    layer1_outputs(6719) <= not(layer0_outputs(8194));
    layer1_outputs(6720) <= not(layer0_outputs(10006));
    layer1_outputs(6721) <= (layer0_outputs(6490)) and (layer0_outputs(10211));
    layer1_outputs(6722) <= layer0_outputs(3778);
    layer1_outputs(6723) <= not((layer0_outputs(4308)) xor (layer0_outputs(4440)));
    layer1_outputs(6724) <= layer0_outputs(3642);
    layer1_outputs(6725) <= not(layer0_outputs(1985));
    layer1_outputs(6726) <= layer0_outputs(5618);
    layer1_outputs(6727) <= (layer0_outputs(9702)) and (layer0_outputs(10058));
    layer1_outputs(6728) <= not((layer0_outputs(6597)) xor (layer0_outputs(8410)));
    layer1_outputs(6729) <= not(layer0_outputs(3169));
    layer1_outputs(6730) <= not((layer0_outputs(1077)) and (layer0_outputs(8812)));
    layer1_outputs(6731) <= not((layer0_outputs(7404)) and (layer0_outputs(1168)));
    layer1_outputs(6732) <= (layer0_outputs(6448)) and (layer0_outputs(107));
    layer1_outputs(6733) <= (layer0_outputs(654)) and (layer0_outputs(7428));
    layer1_outputs(6734) <= (layer0_outputs(1883)) and (layer0_outputs(8451));
    layer1_outputs(6735) <= not(layer0_outputs(7732));
    layer1_outputs(6736) <= not((layer0_outputs(10219)) xor (layer0_outputs(4032)));
    layer1_outputs(6737) <= (layer0_outputs(6810)) or (layer0_outputs(9130));
    layer1_outputs(6738) <= not(layer0_outputs(7553)) or (layer0_outputs(1306));
    layer1_outputs(6739) <= not((layer0_outputs(1104)) or (layer0_outputs(6008)));
    layer1_outputs(6740) <= not((layer0_outputs(5646)) and (layer0_outputs(236)));
    layer1_outputs(6741) <= layer0_outputs(4715);
    layer1_outputs(6742) <= (layer0_outputs(1014)) and (layer0_outputs(3732));
    layer1_outputs(6743) <= not(layer0_outputs(9327));
    layer1_outputs(6744) <= layer0_outputs(916);
    layer1_outputs(6745) <= not(layer0_outputs(9215)) or (layer0_outputs(3708));
    layer1_outputs(6746) <= not(layer0_outputs(1861)) or (layer0_outputs(6348));
    layer1_outputs(6747) <= not(layer0_outputs(1585)) or (layer0_outputs(9749));
    layer1_outputs(6748) <= not((layer0_outputs(1402)) xor (layer0_outputs(1401)));
    layer1_outputs(6749) <= not(layer0_outputs(2748));
    layer1_outputs(6750) <= layer0_outputs(6554);
    layer1_outputs(6751) <= not(layer0_outputs(345)) or (layer0_outputs(559));
    layer1_outputs(6752) <= layer0_outputs(543);
    layer1_outputs(6753) <= (layer0_outputs(2750)) and not (layer0_outputs(6015));
    layer1_outputs(6754) <= not(layer0_outputs(6053));
    layer1_outputs(6755) <= '1';
    layer1_outputs(6756) <= (layer0_outputs(2546)) and (layer0_outputs(9029));
    layer1_outputs(6757) <= not(layer0_outputs(4515));
    layer1_outputs(6758) <= layer0_outputs(2389);
    layer1_outputs(6759) <= '1';
    layer1_outputs(6760) <= (layer0_outputs(1614)) or (layer0_outputs(8497));
    layer1_outputs(6761) <= (layer0_outputs(3935)) and not (layer0_outputs(9358));
    layer1_outputs(6762) <= '1';
    layer1_outputs(6763) <= layer0_outputs(6104);
    layer1_outputs(6764) <= not((layer0_outputs(9855)) or (layer0_outputs(3566)));
    layer1_outputs(6765) <= not(layer0_outputs(8489)) or (layer0_outputs(652));
    layer1_outputs(6766) <= layer0_outputs(6088);
    layer1_outputs(6767) <= (layer0_outputs(6637)) and (layer0_outputs(4938));
    layer1_outputs(6768) <= (layer0_outputs(5889)) and not (layer0_outputs(7545));
    layer1_outputs(6769) <= not(layer0_outputs(6876));
    layer1_outputs(6770) <= not(layer0_outputs(3125));
    layer1_outputs(6771) <= not(layer0_outputs(3942)) or (layer0_outputs(2268));
    layer1_outputs(6772) <= not(layer0_outputs(2641));
    layer1_outputs(6773) <= layer0_outputs(7677);
    layer1_outputs(6774) <= not((layer0_outputs(4168)) xor (layer0_outputs(3067)));
    layer1_outputs(6775) <= not((layer0_outputs(5893)) and (layer0_outputs(6136)));
    layer1_outputs(6776) <= not(layer0_outputs(5985));
    layer1_outputs(6777) <= layer0_outputs(3526);
    layer1_outputs(6778) <= layer0_outputs(7469);
    layer1_outputs(6779) <= not((layer0_outputs(1931)) xor (layer0_outputs(6376)));
    layer1_outputs(6780) <= not((layer0_outputs(6542)) or (layer0_outputs(3504)));
    layer1_outputs(6781) <= layer0_outputs(4043);
    layer1_outputs(6782) <= not(layer0_outputs(597));
    layer1_outputs(6783) <= '0';
    layer1_outputs(6784) <= not(layer0_outputs(8644));
    layer1_outputs(6785) <= layer0_outputs(8379);
    layer1_outputs(6786) <= not(layer0_outputs(7849));
    layer1_outputs(6787) <= not((layer0_outputs(2681)) and (layer0_outputs(4864)));
    layer1_outputs(6788) <= layer0_outputs(1494);
    layer1_outputs(6789) <= layer0_outputs(7451);
    layer1_outputs(6790) <= not((layer0_outputs(5439)) and (layer0_outputs(4746)));
    layer1_outputs(6791) <= not(layer0_outputs(5736));
    layer1_outputs(6792) <= not(layer0_outputs(1311));
    layer1_outputs(6793) <= not(layer0_outputs(7553)) or (layer0_outputs(2038));
    layer1_outputs(6794) <= not((layer0_outputs(8889)) and (layer0_outputs(6055)));
    layer1_outputs(6795) <= (layer0_outputs(7801)) or (layer0_outputs(2041));
    layer1_outputs(6796) <= not(layer0_outputs(10129));
    layer1_outputs(6797) <= '0';
    layer1_outputs(6798) <= '0';
    layer1_outputs(6799) <= (layer0_outputs(2935)) or (layer0_outputs(8620));
    layer1_outputs(6800) <= not(layer0_outputs(1974));
    layer1_outputs(6801) <= (layer0_outputs(10)) and not (layer0_outputs(2992));
    layer1_outputs(6802) <= (layer0_outputs(358)) xor (layer0_outputs(3543));
    layer1_outputs(6803) <= (layer0_outputs(2146)) or (layer0_outputs(7912));
    layer1_outputs(6804) <= not((layer0_outputs(7381)) and (layer0_outputs(2131)));
    layer1_outputs(6805) <= (layer0_outputs(6320)) and not (layer0_outputs(3675));
    layer1_outputs(6806) <= layer0_outputs(7137);
    layer1_outputs(6807) <= layer0_outputs(5924);
    layer1_outputs(6808) <= not((layer0_outputs(8389)) and (layer0_outputs(5460)));
    layer1_outputs(6809) <= layer0_outputs(7939);
    layer1_outputs(6810) <= (layer0_outputs(10083)) and not (layer0_outputs(8116));
    layer1_outputs(6811) <= layer0_outputs(8721);
    layer1_outputs(6812) <= not(layer0_outputs(7116)) or (layer0_outputs(5403));
    layer1_outputs(6813) <= (layer0_outputs(2052)) and (layer0_outputs(171));
    layer1_outputs(6814) <= not(layer0_outputs(2463)) or (layer0_outputs(7757));
    layer1_outputs(6815) <= not(layer0_outputs(5658));
    layer1_outputs(6816) <= (layer0_outputs(5928)) and not (layer0_outputs(153));
    layer1_outputs(6817) <= (layer0_outputs(4274)) and not (layer0_outputs(996));
    layer1_outputs(6818) <= not((layer0_outputs(3455)) or (layer0_outputs(4489)));
    layer1_outputs(6819) <= not(layer0_outputs(8308));
    layer1_outputs(6820) <= not((layer0_outputs(6758)) or (layer0_outputs(9659)));
    layer1_outputs(6821) <= not(layer0_outputs(0));
    layer1_outputs(6822) <= (layer0_outputs(9369)) or (layer0_outputs(6720));
    layer1_outputs(6823) <= (layer0_outputs(10086)) or (layer0_outputs(5523));
    layer1_outputs(6824) <= not((layer0_outputs(5600)) and (layer0_outputs(1333)));
    layer1_outputs(6825) <= (layer0_outputs(7020)) and not (layer0_outputs(6291));
    layer1_outputs(6826) <= (layer0_outputs(2110)) and not (layer0_outputs(6195));
    layer1_outputs(6827) <= not(layer0_outputs(4385)) or (layer0_outputs(4974));
    layer1_outputs(6828) <= (layer0_outputs(7623)) xor (layer0_outputs(3268));
    layer1_outputs(6829) <= not(layer0_outputs(805));
    layer1_outputs(6830) <= (layer0_outputs(6408)) and (layer0_outputs(5989));
    layer1_outputs(6831) <= not(layer0_outputs(353));
    layer1_outputs(6832) <= not(layer0_outputs(5992));
    layer1_outputs(6833) <= not((layer0_outputs(1721)) and (layer0_outputs(8899)));
    layer1_outputs(6834) <= not(layer0_outputs(4544));
    layer1_outputs(6835) <= not((layer0_outputs(5337)) xor (layer0_outputs(558)));
    layer1_outputs(6836) <= (layer0_outputs(5605)) xor (layer0_outputs(6036));
    layer1_outputs(6837) <= (layer0_outputs(2025)) or (layer0_outputs(829));
    layer1_outputs(6838) <= not(layer0_outputs(4265));
    layer1_outputs(6839) <= not((layer0_outputs(8372)) or (layer0_outputs(3828)));
    layer1_outputs(6840) <= not(layer0_outputs(3735));
    layer1_outputs(6841) <= layer0_outputs(9135);
    layer1_outputs(6842) <= not(layer0_outputs(5140));
    layer1_outputs(6843) <= not(layer0_outputs(2085)) or (layer0_outputs(3850));
    layer1_outputs(6844) <= layer0_outputs(8506);
    layer1_outputs(6845) <= not(layer0_outputs(5723));
    layer1_outputs(6846) <= not(layer0_outputs(5792)) or (layer0_outputs(9774));
    layer1_outputs(6847) <= not(layer0_outputs(7119));
    layer1_outputs(6848) <= layer0_outputs(1499);
    layer1_outputs(6849) <= not(layer0_outputs(5699));
    layer1_outputs(6850) <= (layer0_outputs(1357)) or (layer0_outputs(6390));
    layer1_outputs(6851) <= not(layer0_outputs(9435));
    layer1_outputs(6852) <= (layer0_outputs(4618)) and not (layer0_outputs(6227));
    layer1_outputs(6853) <= (layer0_outputs(1859)) and not (layer0_outputs(136));
    layer1_outputs(6854) <= not((layer0_outputs(5432)) xor (layer0_outputs(2810)));
    layer1_outputs(6855) <= (layer0_outputs(2798)) and not (layer0_outputs(418));
    layer1_outputs(6856) <= not((layer0_outputs(7126)) xor (layer0_outputs(686)));
    layer1_outputs(6857) <= not(layer0_outputs(784));
    layer1_outputs(6858) <= not((layer0_outputs(798)) or (layer0_outputs(5429)));
    layer1_outputs(6859) <= layer0_outputs(4979);
    layer1_outputs(6860) <= not(layer0_outputs(9868)) or (layer0_outputs(5270));
    layer1_outputs(6861) <= layer0_outputs(7268);
    layer1_outputs(6862) <= (layer0_outputs(6845)) or (layer0_outputs(2631));
    layer1_outputs(6863) <= not((layer0_outputs(7850)) and (layer0_outputs(2092)));
    layer1_outputs(6864) <= not((layer0_outputs(611)) xor (layer0_outputs(7898)));
    layer1_outputs(6865) <= not(layer0_outputs(9343));
    layer1_outputs(6866) <= layer0_outputs(8330);
    layer1_outputs(6867) <= not(layer0_outputs(9097)) or (layer0_outputs(5112));
    layer1_outputs(6868) <= layer0_outputs(5022);
    layer1_outputs(6869) <= not((layer0_outputs(1903)) and (layer0_outputs(2573)));
    layer1_outputs(6870) <= not(layer0_outputs(5746)) or (layer0_outputs(2762));
    layer1_outputs(6871) <= not((layer0_outputs(2494)) and (layer0_outputs(2619)));
    layer1_outputs(6872) <= layer0_outputs(6781);
    layer1_outputs(6873) <= (layer0_outputs(7675)) and not (layer0_outputs(161));
    layer1_outputs(6874) <= (layer0_outputs(5965)) and (layer0_outputs(3714));
    layer1_outputs(6875) <= (layer0_outputs(5631)) and not (layer0_outputs(2724));
    layer1_outputs(6876) <= (layer0_outputs(2647)) and not (layer0_outputs(7533));
    layer1_outputs(6877) <= (layer0_outputs(7510)) and not (layer0_outputs(9212));
    layer1_outputs(6878) <= layer0_outputs(2227);
    layer1_outputs(6879) <= layer0_outputs(1584);
    layer1_outputs(6880) <= layer0_outputs(8088);
    layer1_outputs(6881) <= not((layer0_outputs(8893)) and (layer0_outputs(6144)));
    layer1_outputs(6882) <= not(layer0_outputs(7894));
    layer1_outputs(6883) <= (layer0_outputs(6807)) and not (layer0_outputs(863));
    layer1_outputs(6884) <= '0';
    layer1_outputs(6885) <= (layer0_outputs(5685)) and not (layer0_outputs(7259));
    layer1_outputs(6886) <= layer0_outputs(6775);
    layer1_outputs(6887) <= not((layer0_outputs(3235)) or (layer0_outputs(8020)));
    layer1_outputs(6888) <= not(layer0_outputs(4465));
    layer1_outputs(6889) <= not((layer0_outputs(8492)) and (layer0_outputs(9037)));
    layer1_outputs(6890) <= not((layer0_outputs(4261)) xor (layer0_outputs(459)));
    layer1_outputs(6891) <= layer0_outputs(5947);
    layer1_outputs(6892) <= not((layer0_outputs(9787)) or (layer0_outputs(7855)));
    layer1_outputs(6893) <= (layer0_outputs(7960)) and not (layer0_outputs(2241));
    layer1_outputs(6894) <= not(layer0_outputs(4154));
    layer1_outputs(6895) <= layer0_outputs(6160);
    layer1_outputs(6896) <= not((layer0_outputs(4912)) and (layer0_outputs(7999)));
    layer1_outputs(6897) <= not(layer0_outputs(369));
    layer1_outputs(6898) <= (layer0_outputs(9608)) or (layer0_outputs(5328));
    layer1_outputs(6899) <= (layer0_outputs(9677)) and not (layer0_outputs(5274));
    layer1_outputs(6900) <= not(layer0_outputs(1569));
    layer1_outputs(6901) <= not((layer0_outputs(6022)) xor (layer0_outputs(5751)));
    layer1_outputs(6902) <= (layer0_outputs(10002)) xor (layer0_outputs(922));
    layer1_outputs(6903) <= not(layer0_outputs(9886));
    layer1_outputs(6904) <= layer0_outputs(6600);
    layer1_outputs(6905) <= layer0_outputs(7861);
    layer1_outputs(6906) <= not(layer0_outputs(8384)) or (layer0_outputs(5804));
    layer1_outputs(6907) <= not(layer0_outputs(1696));
    layer1_outputs(6908) <= '1';
    layer1_outputs(6909) <= layer0_outputs(1131);
    layer1_outputs(6910) <= (layer0_outputs(3412)) and not (layer0_outputs(826));
    layer1_outputs(6911) <= not(layer0_outputs(8049)) or (layer0_outputs(6605));
    layer1_outputs(6912) <= layer0_outputs(3003);
    layer1_outputs(6913) <= '0';
    layer1_outputs(6914) <= (layer0_outputs(17)) or (layer0_outputs(9273));
    layer1_outputs(6915) <= (layer0_outputs(9763)) and not (layer0_outputs(2261));
    layer1_outputs(6916) <= not(layer0_outputs(4157));
    layer1_outputs(6917) <= not(layer0_outputs(2621)) or (layer0_outputs(1300));
    layer1_outputs(6918) <= not(layer0_outputs(2783));
    layer1_outputs(6919) <= not((layer0_outputs(2928)) or (layer0_outputs(7062)));
    layer1_outputs(6920) <= layer0_outputs(1382);
    layer1_outputs(6921) <= not(layer0_outputs(579));
    layer1_outputs(6922) <= (layer0_outputs(4008)) or (layer0_outputs(4582));
    layer1_outputs(6923) <= layer0_outputs(6340);
    layer1_outputs(6924) <= layer0_outputs(8728);
    layer1_outputs(6925) <= not((layer0_outputs(9289)) and (layer0_outputs(9476)));
    layer1_outputs(6926) <= not(layer0_outputs(1985)) or (layer0_outputs(9679));
    layer1_outputs(6927) <= (layer0_outputs(5177)) and not (layer0_outputs(9541));
    layer1_outputs(6928) <= (layer0_outputs(118)) and not (layer0_outputs(6351));
    layer1_outputs(6929) <= layer0_outputs(8627);
    layer1_outputs(6930) <= (layer0_outputs(8375)) or (layer0_outputs(6952));
    layer1_outputs(6931) <= not((layer0_outputs(3884)) or (layer0_outputs(9090)));
    layer1_outputs(6932) <= layer0_outputs(4660);
    layer1_outputs(6933) <= not(layer0_outputs(687));
    layer1_outputs(6934) <= layer0_outputs(4804);
    layer1_outputs(6935) <= not(layer0_outputs(6827));
    layer1_outputs(6936) <= (layer0_outputs(1500)) and (layer0_outputs(2409));
    layer1_outputs(6937) <= not((layer0_outputs(2111)) or (layer0_outputs(3015)));
    layer1_outputs(6938) <= not(layer0_outputs(4383)) or (layer0_outputs(7324));
    layer1_outputs(6939) <= not(layer0_outputs(5371));
    layer1_outputs(6940) <= (layer0_outputs(563)) or (layer0_outputs(6779));
    layer1_outputs(6941) <= not(layer0_outputs(4823)) or (layer0_outputs(3878));
    layer1_outputs(6942) <= not(layer0_outputs(2435));
    layer1_outputs(6943) <= (layer0_outputs(8466)) xor (layer0_outputs(2243));
    layer1_outputs(6944) <= not((layer0_outputs(9087)) and (layer0_outputs(7499)));
    layer1_outputs(6945) <= not((layer0_outputs(5161)) xor (layer0_outputs(2286)));
    layer1_outputs(6946) <= not(layer0_outputs(3683));
    layer1_outputs(6947) <= layer0_outputs(2781);
    layer1_outputs(6948) <= not((layer0_outputs(1866)) or (layer0_outputs(3069)));
    layer1_outputs(6949) <= not(layer0_outputs(3904));
    layer1_outputs(6950) <= not((layer0_outputs(7073)) and (layer0_outputs(644)));
    layer1_outputs(6951) <= not(layer0_outputs(8244));
    layer1_outputs(6952) <= (layer0_outputs(2367)) and not (layer0_outputs(2146));
    layer1_outputs(6953) <= not(layer0_outputs(2792)) or (layer0_outputs(7874));
    layer1_outputs(6954) <= layer0_outputs(9736);
    layer1_outputs(6955) <= layer0_outputs(9866);
    layer1_outputs(6956) <= not(layer0_outputs(1572)) or (layer0_outputs(10175));
    layer1_outputs(6957) <= not((layer0_outputs(182)) and (layer0_outputs(9460)));
    layer1_outputs(6958) <= not(layer0_outputs(4655)) or (layer0_outputs(10157));
    layer1_outputs(6959) <= not((layer0_outputs(6568)) and (layer0_outputs(8211)));
    layer1_outputs(6960) <= not((layer0_outputs(3527)) or (layer0_outputs(4769)));
    layer1_outputs(6961) <= layer0_outputs(8109);
    layer1_outputs(6962) <= layer0_outputs(8129);
    layer1_outputs(6963) <= layer0_outputs(2615);
    layer1_outputs(6964) <= '0';
    layer1_outputs(6965) <= not(layer0_outputs(9462)) or (layer0_outputs(4499));
    layer1_outputs(6966) <= (layer0_outputs(4424)) and not (layer0_outputs(6980));
    layer1_outputs(6967) <= not(layer0_outputs(9531));
    layer1_outputs(6968) <= not(layer0_outputs(2901));
    layer1_outputs(6969) <= not(layer0_outputs(3625)) or (layer0_outputs(6534));
    layer1_outputs(6970) <= layer0_outputs(1998);
    layer1_outputs(6971) <= (layer0_outputs(3827)) or (layer0_outputs(2353));
    layer1_outputs(6972) <= not(layer0_outputs(8572));
    layer1_outputs(6973) <= layer0_outputs(6572);
    layer1_outputs(6974) <= layer0_outputs(7724);
    layer1_outputs(6975) <= layer0_outputs(7942);
    layer1_outputs(6976) <= not(layer0_outputs(1901));
    layer1_outputs(6977) <= (layer0_outputs(8578)) and (layer0_outputs(8596));
    layer1_outputs(6978) <= not(layer0_outputs(3298)) or (layer0_outputs(3479));
    layer1_outputs(6979) <= layer0_outputs(6337);
    layer1_outputs(6980) <= layer0_outputs(3424);
    layer1_outputs(6981) <= not(layer0_outputs(8595));
    layer1_outputs(6982) <= (layer0_outputs(9153)) and (layer0_outputs(1474));
    layer1_outputs(6983) <= not((layer0_outputs(1172)) or (layer0_outputs(10212)));
    layer1_outputs(6984) <= layer0_outputs(8260);
    layer1_outputs(6985) <= (layer0_outputs(4393)) or (layer0_outputs(6621));
    layer1_outputs(6986) <= not((layer0_outputs(5653)) and (layer0_outputs(7177)));
    layer1_outputs(6987) <= not((layer0_outputs(5597)) or (layer0_outputs(4493)));
    layer1_outputs(6988) <= '0';
    layer1_outputs(6989) <= (layer0_outputs(3328)) and (layer0_outputs(7668));
    layer1_outputs(6990) <= (layer0_outputs(4587)) and not (layer0_outputs(5247));
    layer1_outputs(6991) <= '1';
    layer1_outputs(6992) <= layer0_outputs(3629);
    layer1_outputs(6993) <= (layer0_outputs(6993)) and (layer0_outputs(8510));
    layer1_outputs(6994) <= not((layer0_outputs(3442)) or (layer0_outputs(6602)));
    layer1_outputs(6995) <= (layer0_outputs(4761)) or (layer0_outputs(8158));
    layer1_outputs(6996) <= not(layer0_outputs(10098)) or (layer0_outputs(1355));
    layer1_outputs(6997) <= layer0_outputs(639);
    layer1_outputs(6998) <= (layer0_outputs(8451)) xor (layer0_outputs(6065));
    layer1_outputs(6999) <= not(layer0_outputs(9782));
    layer1_outputs(7000) <= (layer0_outputs(9169)) and not (layer0_outputs(6752));
    layer1_outputs(7001) <= layer0_outputs(1201);
    layer1_outputs(7002) <= layer0_outputs(5358);
    layer1_outputs(7003) <= (layer0_outputs(1982)) and not (layer0_outputs(5116));
    layer1_outputs(7004) <= layer0_outputs(6121);
    layer1_outputs(7005) <= (layer0_outputs(413)) xor (layer0_outputs(9112));
    layer1_outputs(7006) <= (layer0_outputs(742)) and not (layer0_outputs(9075));
    layer1_outputs(7007) <= not(layer0_outputs(1370));
    layer1_outputs(7008) <= not(layer0_outputs(1223)) or (layer0_outputs(9996));
    layer1_outputs(7009) <= (layer0_outputs(3666)) or (layer0_outputs(227));
    layer1_outputs(7010) <= not((layer0_outputs(7735)) and (layer0_outputs(640)));
    layer1_outputs(7011) <= layer0_outputs(9105);
    layer1_outputs(7012) <= not((layer0_outputs(5945)) or (layer0_outputs(4097)));
    layer1_outputs(7013) <= layer0_outputs(9793);
    layer1_outputs(7014) <= (layer0_outputs(6398)) xor (layer0_outputs(6016));
    layer1_outputs(7015) <= (layer0_outputs(474)) xor (layer0_outputs(9937));
    layer1_outputs(7016) <= not(layer0_outputs(9314));
    layer1_outputs(7017) <= (layer0_outputs(5498)) xor (layer0_outputs(734));
    layer1_outputs(7018) <= layer0_outputs(6879);
    layer1_outputs(7019) <= not(layer0_outputs(8969));
    layer1_outputs(7020) <= (layer0_outputs(5130)) or (layer0_outputs(4108));
    layer1_outputs(7021) <= not(layer0_outputs(912)) or (layer0_outputs(7357));
    layer1_outputs(7022) <= not(layer0_outputs(2167));
    layer1_outputs(7023) <= not(layer0_outputs(5784)) or (layer0_outputs(2462));
    layer1_outputs(7024) <= (layer0_outputs(7046)) xor (layer0_outputs(3041));
    layer1_outputs(7025) <= not(layer0_outputs(2272));
    layer1_outputs(7026) <= not(layer0_outputs(6538));
    layer1_outputs(7027) <= layer0_outputs(2822);
    layer1_outputs(7028) <= not(layer0_outputs(9596));
    layer1_outputs(7029) <= not(layer0_outputs(9711));
    layer1_outputs(7030) <= layer0_outputs(7728);
    layer1_outputs(7031) <= (layer0_outputs(5696)) or (layer0_outputs(3902));
    layer1_outputs(7032) <= layer0_outputs(7984);
    layer1_outputs(7033) <= layer0_outputs(5144);
    layer1_outputs(7034) <= not(layer0_outputs(10042)) or (layer0_outputs(2320));
    layer1_outputs(7035) <= not((layer0_outputs(8376)) xor (layer0_outputs(2047)));
    layer1_outputs(7036) <= not(layer0_outputs(6208));
    layer1_outputs(7037) <= layer0_outputs(1855);
    layer1_outputs(7038) <= (layer0_outputs(2133)) xor (layer0_outputs(7720));
    layer1_outputs(7039) <= (layer0_outputs(1258)) and (layer0_outputs(999));
    layer1_outputs(7040) <= not((layer0_outputs(7248)) and (layer0_outputs(4952)));
    layer1_outputs(7041) <= (layer0_outputs(7905)) xor (layer0_outputs(1758));
    layer1_outputs(7042) <= not(layer0_outputs(6256));
    layer1_outputs(7043) <= layer0_outputs(8169);
    layer1_outputs(7044) <= (layer0_outputs(9479)) and not (layer0_outputs(8125));
    layer1_outputs(7045) <= not((layer0_outputs(9929)) or (layer0_outputs(1910)));
    layer1_outputs(7046) <= not(layer0_outputs(6064));
    layer1_outputs(7047) <= layer0_outputs(5956);
    layer1_outputs(7048) <= not(layer0_outputs(4250)) or (layer0_outputs(1193));
    layer1_outputs(7049) <= layer0_outputs(5142);
    layer1_outputs(7050) <= not(layer0_outputs(9259));
    layer1_outputs(7051) <= (layer0_outputs(5238)) and not (layer0_outputs(4574));
    layer1_outputs(7052) <= '1';
    layer1_outputs(7053) <= layer0_outputs(68);
    layer1_outputs(7054) <= not(layer0_outputs(7130)) or (layer0_outputs(3200));
    layer1_outputs(7055) <= not(layer0_outputs(1146));
    layer1_outputs(7056) <= not(layer0_outputs(3794));
    layer1_outputs(7057) <= not(layer0_outputs(2508));
    layer1_outputs(7058) <= not(layer0_outputs(1338));
    layer1_outputs(7059) <= (layer0_outputs(10070)) and not (layer0_outputs(6102));
    layer1_outputs(7060) <= (layer0_outputs(1024)) and (layer0_outputs(5445));
    layer1_outputs(7061) <= (layer0_outputs(4968)) and (layer0_outputs(7140));
    layer1_outputs(7062) <= (layer0_outputs(3063)) or (layer0_outputs(7580));
    layer1_outputs(7063) <= not(layer0_outputs(4049));
    layer1_outputs(7064) <= (layer0_outputs(8120)) and not (layer0_outputs(2836));
    layer1_outputs(7065) <= not(layer0_outputs(9432)) or (layer0_outputs(4515));
    layer1_outputs(7066) <= not(layer0_outputs(8044));
    layer1_outputs(7067) <= not(layer0_outputs(6652));
    layer1_outputs(7068) <= '0';
    layer1_outputs(7069) <= not(layer0_outputs(2670));
    layer1_outputs(7070) <= layer0_outputs(6143);
    layer1_outputs(7071) <= '0';
    layer1_outputs(7072) <= not((layer0_outputs(2540)) xor (layer0_outputs(5588)));
    layer1_outputs(7073) <= not(layer0_outputs(30));
    layer1_outputs(7074) <= layer0_outputs(1682);
    layer1_outputs(7075) <= (layer0_outputs(5979)) and not (layer0_outputs(10101));
    layer1_outputs(7076) <= (layer0_outputs(2530)) or (layer0_outputs(2824));
    layer1_outputs(7077) <= '0';
    layer1_outputs(7078) <= not(layer0_outputs(9574)) or (layer0_outputs(9879));
    layer1_outputs(7079) <= layer0_outputs(3757);
    layer1_outputs(7080) <= not((layer0_outputs(2350)) or (layer0_outputs(8670)));
    layer1_outputs(7081) <= (layer0_outputs(4394)) and not (layer0_outputs(9816));
    layer1_outputs(7082) <= '1';
    layer1_outputs(7083) <= '0';
    layer1_outputs(7084) <= (layer0_outputs(6248)) and (layer0_outputs(4260));
    layer1_outputs(7085) <= layer0_outputs(2888);
    layer1_outputs(7086) <= '0';
    layer1_outputs(7087) <= (layer0_outputs(8757)) xor (layer0_outputs(882));
    layer1_outputs(7088) <= (layer0_outputs(9487)) and not (layer0_outputs(6917));
    layer1_outputs(7089) <= not(layer0_outputs(1378));
    layer1_outputs(7090) <= not(layer0_outputs(1307));
    layer1_outputs(7091) <= layer0_outputs(5629);
    layer1_outputs(7092) <= not(layer0_outputs(6250));
    layer1_outputs(7093) <= not(layer0_outputs(9145));
    layer1_outputs(7094) <= not(layer0_outputs(8828)) or (layer0_outputs(1181));
    layer1_outputs(7095) <= (layer0_outputs(8024)) or (layer0_outputs(1419));
    layer1_outputs(7096) <= not(layer0_outputs(3787));
    layer1_outputs(7097) <= '1';
    layer1_outputs(7098) <= not(layer0_outputs(6200)) or (layer0_outputs(335));
    layer1_outputs(7099) <= not((layer0_outputs(3591)) or (layer0_outputs(9903)));
    layer1_outputs(7100) <= not((layer0_outputs(3032)) or (layer0_outputs(5940)));
    layer1_outputs(7101) <= (layer0_outputs(6494)) or (layer0_outputs(10144));
    layer1_outputs(7102) <= not((layer0_outputs(7607)) or (layer0_outputs(7767)));
    layer1_outputs(7103) <= layer0_outputs(1233);
    layer1_outputs(7104) <= not((layer0_outputs(3907)) xor (layer0_outputs(4534)));
    layer1_outputs(7105) <= (layer0_outputs(7959)) or (layer0_outputs(1884));
    layer1_outputs(7106) <= not(layer0_outputs(1595));
    layer1_outputs(7107) <= not((layer0_outputs(5168)) and (layer0_outputs(4565)));
    layer1_outputs(7108) <= layer0_outputs(3155);
    layer1_outputs(7109) <= (layer0_outputs(5690)) and (layer0_outputs(6530));
    layer1_outputs(7110) <= not(layer0_outputs(5708));
    layer1_outputs(7111) <= layer0_outputs(123);
    layer1_outputs(7112) <= (layer0_outputs(8218)) and (layer0_outputs(2264));
    layer1_outputs(7113) <= not(layer0_outputs(3030));
    layer1_outputs(7114) <= not((layer0_outputs(207)) or (layer0_outputs(7917)));
    layer1_outputs(7115) <= layer0_outputs(1788);
    layer1_outputs(7116) <= (layer0_outputs(9134)) and not (layer0_outputs(7830));
    layer1_outputs(7117) <= not((layer0_outputs(8071)) xor (layer0_outputs(7039)));
    layer1_outputs(7118) <= not(layer0_outputs(2988));
    layer1_outputs(7119) <= layer0_outputs(5126);
    layer1_outputs(7120) <= not(layer0_outputs(7038));
    layer1_outputs(7121) <= not(layer0_outputs(1078)) or (layer0_outputs(3511));
    layer1_outputs(7122) <= layer0_outputs(9185);
    layer1_outputs(7123) <= not(layer0_outputs(7695)) or (layer0_outputs(7569));
    layer1_outputs(7124) <= (layer0_outputs(2666)) and (layer0_outputs(3839));
    layer1_outputs(7125) <= not(layer0_outputs(6976));
    layer1_outputs(7126) <= (layer0_outputs(6804)) and not (layer0_outputs(5649));
    layer1_outputs(7127) <= not(layer0_outputs(3258));
    layer1_outputs(7128) <= '1';
    layer1_outputs(7129) <= not(layer0_outputs(4058));
    layer1_outputs(7130) <= not(layer0_outputs(4079));
    layer1_outputs(7131) <= layer0_outputs(2104);
    layer1_outputs(7132) <= (layer0_outputs(5036)) and (layer0_outputs(3418));
    layer1_outputs(7133) <= not((layer0_outputs(656)) and (layer0_outputs(6302)));
    layer1_outputs(7134) <= not(layer0_outputs(3585)) or (layer0_outputs(4079));
    layer1_outputs(7135) <= not(layer0_outputs(2999));
    layer1_outputs(7136) <= not((layer0_outputs(6861)) xor (layer0_outputs(3564)));
    layer1_outputs(7137) <= (layer0_outputs(7344)) and not (layer0_outputs(8973));
    layer1_outputs(7138) <= not(layer0_outputs(2397)) or (layer0_outputs(5169));
    layer1_outputs(7139) <= not(layer0_outputs(2308)) or (layer0_outputs(4461));
    layer1_outputs(7140) <= '0';
    layer1_outputs(7141) <= (layer0_outputs(4111)) and (layer0_outputs(7749));
    layer1_outputs(7142) <= not((layer0_outputs(3666)) and (layer0_outputs(9502)));
    layer1_outputs(7143) <= not(layer0_outputs(3019)) or (layer0_outputs(6067));
    layer1_outputs(7144) <= not((layer0_outputs(3769)) and (layer0_outputs(8859)));
    layer1_outputs(7145) <= not(layer0_outputs(8620));
    layer1_outputs(7146) <= (layer0_outputs(8845)) and not (layer0_outputs(4712));
    layer1_outputs(7147) <= '0';
    layer1_outputs(7148) <= not((layer0_outputs(9938)) and (layer0_outputs(7185)));
    layer1_outputs(7149) <= not(layer0_outputs(7389));
    layer1_outputs(7150) <= (layer0_outputs(8880)) and not (layer0_outputs(6219));
    layer1_outputs(7151) <= not((layer0_outputs(6675)) or (layer0_outputs(3097)));
    layer1_outputs(7152) <= (layer0_outputs(8277)) and (layer0_outputs(3667));
    layer1_outputs(7153) <= not((layer0_outputs(3582)) and (layer0_outputs(9155)));
    layer1_outputs(7154) <= not(layer0_outputs(3052)) or (layer0_outputs(5824));
    layer1_outputs(7155) <= (layer0_outputs(4816)) and not (layer0_outputs(188));
    layer1_outputs(7156) <= not((layer0_outputs(3232)) xor (layer0_outputs(423)));
    layer1_outputs(7157) <= not((layer0_outputs(1094)) and (layer0_outputs(6137)));
    layer1_outputs(7158) <= (layer0_outputs(3263)) or (layer0_outputs(3749));
    layer1_outputs(7159) <= layer0_outputs(5030);
    layer1_outputs(7160) <= not((layer0_outputs(7966)) or (layer0_outputs(1139)));
    layer1_outputs(7161) <= layer0_outputs(2150);
    layer1_outputs(7162) <= not(layer0_outputs(528));
    layer1_outputs(7163) <= layer0_outputs(9624);
    layer1_outputs(7164) <= not((layer0_outputs(4744)) or (layer0_outputs(5324)));
    layer1_outputs(7165) <= not(layer0_outputs(1583));
    layer1_outputs(7166) <= (layer0_outputs(7994)) or (layer0_outputs(1454));
    layer1_outputs(7167) <= (layer0_outputs(3347)) and not (layer0_outputs(7945));
    layer1_outputs(7168) <= layer0_outputs(8156);
    layer1_outputs(7169) <= (layer0_outputs(8624)) and not (layer0_outputs(738));
    layer1_outputs(7170) <= not((layer0_outputs(2386)) and (layer0_outputs(7682)));
    layer1_outputs(7171) <= not((layer0_outputs(3072)) or (layer0_outputs(7419)));
    layer1_outputs(7172) <= not(layer0_outputs(8739));
    layer1_outputs(7173) <= layer0_outputs(5210);
    layer1_outputs(7174) <= not(layer0_outputs(551));
    layer1_outputs(7175) <= not((layer0_outputs(6920)) or (layer0_outputs(8453)));
    layer1_outputs(7176) <= not(layer0_outputs(700)) or (layer0_outputs(2053));
    layer1_outputs(7177) <= not(layer0_outputs(880));
    layer1_outputs(7178) <= (layer0_outputs(6400)) and not (layer0_outputs(5175));
    layer1_outputs(7179) <= not(layer0_outputs(627)) or (layer0_outputs(2949));
    layer1_outputs(7180) <= not(layer0_outputs(7364)) or (layer0_outputs(5264));
    layer1_outputs(7181) <= not((layer0_outputs(7330)) xor (layer0_outputs(5737)));
    layer1_outputs(7182) <= layer0_outputs(6749);
    layer1_outputs(7183) <= (layer0_outputs(8332)) or (layer0_outputs(7029));
    layer1_outputs(7184) <= layer0_outputs(8685);
    layer1_outputs(7185) <= not((layer0_outputs(5537)) xor (layer0_outputs(4007)));
    layer1_outputs(7186) <= not(layer0_outputs(7234)) or (layer0_outputs(9707));
    layer1_outputs(7187) <= not(layer0_outputs(543)) or (layer0_outputs(10194));
    layer1_outputs(7188) <= not(layer0_outputs(8347)) or (layer0_outputs(8462));
    layer1_outputs(7189) <= (layer0_outputs(7620)) xor (layer0_outputs(406));
    layer1_outputs(7190) <= not(layer0_outputs(8633));
    layer1_outputs(7191) <= layer0_outputs(3336);
    layer1_outputs(7192) <= not(layer0_outputs(8585));
    layer1_outputs(7193) <= (layer0_outputs(5007)) and not (layer0_outputs(10011));
    layer1_outputs(7194) <= '0';
    layer1_outputs(7195) <= not(layer0_outputs(8067));
    layer1_outputs(7196) <= '0';
    layer1_outputs(7197) <= not(layer0_outputs(6879));
    layer1_outputs(7198) <= not((layer0_outputs(731)) or (layer0_outputs(4791)));
    layer1_outputs(7199) <= layer0_outputs(4871);
    layer1_outputs(7200) <= (layer0_outputs(7940)) and (layer0_outputs(1673));
    layer1_outputs(7201) <= '1';
    layer1_outputs(7202) <= not(layer0_outputs(5894));
    layer1_outputs(7203) <= not((layer0_outputs(447)) or (layer0_outputs(4361)));
    layer1_outputs(7204) <= (layer0_outputs(4131)) xor (layer0_outputs(7866));
    layer1_outputs(7205) <= not(layer0_outputs(8589));
    layer1_outputs(7206) <= '0';
    layer1_outputs(7207) <= not(layer0_outputs(4528));
    layer1_outputs(7208) <= layer0_outputs(2782);
    layer1_outputs(7209) <= (layer0_outputs(6521)) and not (layer0_outputs(5362));
    layer1_outputs(7210) <= layer0_outputs(8349);
    layer1_outputs(7211) <= (layer0_outputs(3038)) and not (layer0_outputs(4371));
    layer1_outputs(7212) <= not((layer0_outputs(9500)) and (layer0_outputs(7262)));
    layer1_outputs(7213) <= (layer0_outputs(7074)) xor (layer0_outputs(5748));
    layer1_outputs(7214) <= layer0_outputs(2077);
    layer1_outputs(7215) <= '0';
    layer1_outputs(7216) <= not((layer0_outputs(4860)) or (layer0_outputs(307)));
    layer1_outputs(7217) <= not(layer0_outputs(3744)) or (layer0_outputs(4619));
    layer1_outputs(7218) <= not((layer0_outputs(10)) and (layer0_outputs(1277)));
    layer1_outputs(7219) <= layer0_outputs(4695);
    layer1_outputs(7220) <= (layer0_outputs(410)) and not (layer0_outputs(7208));
    layer1_outputs(7221) <= not((layer0_outputs(2312)) and (layer0_outputs(8517)));
    layer1_outputs(7222) <= layer0_outputs(7495);
    layer1_outputs(7223) <= not((layer0_outputs(4395)) or (layer0_outputs(7514)));
    layer1_outputs(7224) <= not((layer0_outputs(6301)) and (layer0_outputs(3739)));
    layer1_outputs(7225) <= not(layer0_outputs(5410)) or (layer0_outputs(8415));
    layer1_outputs(7226) <= layer0_outputs(4426);
    layer1_outputs(7227) <= layer0_outputs(5636);
    layer1_outputs(7228) <= not(layer0_outputs(10126));
    layer1_outputs(7229) <= layer0_outputs(803);
    layer1_outputs(7230) <= (layer0_outputs(3316)) and (layer0_outputs(5378));
    layer1_outputs(7231) <= '1';
    layer1_outputs(7232) <= layer0_outputs(9909);
    layer1_outputs(7233) <= not(layer0_outputs(3017)) or (layer0_outputs(2423));
    layer1_outputs(7234) <= (layer0_outputs(8560)) and not (layer0_outputs(1541));
    layer1_outputs(7235) <= not((layer0_outputs(8241)) and (layer0_outputs(2115)));
    layer1_outputs(7236) <= not(layer0_outputs(8124));
    layer1_outputs(7237) <= layer0_outputs(2411);
    layer1_outputs(7238) <= (layer0_outputs(10085)) or (layer0_outputs(3207));
    layer1_outputs(7239) <= layer0_outputs(6935);
    layer1_outputs(7240) <= layer0_outputs(5708);
    layer1_outputs(7241) <= layer0_outputs(5499);
    layer1_outputs(7242) <= not(layer0_outputs(6096)) or (layer0_outputs(9122));
    layer1_outputs(7243) <= not(layer0_outputs(6650));
    layer1_outputs(7244) <= not(layer0_outputs(6270)) or (layer0_outputs(8965));
    layer1_outputs(7245) <= not(layer0_outputs(10038));
    layer1_outputs(7246) <= not((layer0_outputs(6269)) xor (layer0_outputs(3712)));
    layer1_outputs(7247) <= layer0_outputs(172);
    layer1_outputs(7248) <= not(layer0_outputs(4695));
    layer1_outputs(7249) <= (layer0_outputs(5855)) or (layer0_outputs(8045));
    layer1_outputs(7250) <= (layer0_outputs(2023)) and not (layer0_outputs(5513));
    layer1_outputs(7251) <= not(layer0_outputs(10002)) or (layer0_outputs(9072));
    layer1_outputs(7252) <= layer0_outputs(7850);
    layer1_outputs(7253) <= (layer0_outputs(8735)) and not (layer0_outputs(8906));
    layer1_outputs(7254) <= not(layer0_outputs(52)) or (layer0_outputs(2690));
    layer1_outputs(7255) <= not((layer0_outputs(448)) and (layer0_outputs(671)));
    layer1_outputs(7256) <= layer0_outputs(1275);
    layer1_outputs(7257) <= layer0_outputs(5008);
    layer1_outputs(7258) <= not(layer0_outputs(4813)) or (layer0_outputs(5268));
    layer1_outputs(7259) <= (layer0_outputs(7832)) and not (layer0_outputs(6851));
    layer1_outputs(7260) <= not((layer0_outputs(7182)) and (layer0_outputs(8013)));
    layer1_outputs(7261) <= (layer0_outputs(5860)) xor (layer0_outputs(9811));
    layer1_outputs(7262) <= not(layer0_outputs(9260)) or (layer0_outputs(1397));
    layer1_outputs(7263) <= '1';
    layer1_outputs(7264) <= not(layer0_outputs(2564)) or (layer0_outputs(8656));
    layer1_outputs(7265) <= layer0_outputs(6041);
    layer1_outputs(7266) <= not(layer0_outputs(3409));
    layer1_outputs(7267) <= not(layer0_outputs(6765));
    layer1_outputs(7268) <= layer0_outputs(7931);
    layer1_outputs(7269) <= layer0_outputs(8486);
    layer1_outputs(7270) <= not((layer0_outputs(6214)) xor (layer0_outputs(5998)));
    layer1_outputs(7271) <= (layer0_outputs(8426)) and (layer0_outputs(6819));
    layer1_outputs(7272) <= not((layer0_outputs(6837)) xor (layer0_outputs(3704)));
    layer1_outputs(7273) <= not(layer0_outputs(9983));
    layer1_outputs(7274) <= (layer0_outputs(7893)) and not (layer0_outputs(4442));
    layer1_outputs(7275) <= layer0_outputs(7978);
    layer1_outputs(7276) <= (layer0_outputs(604)) and not (layer0_outputs(2978));
    layer1_outputs(7277) <= '0';
    layer1_outputs(7278) <= not((layer0_outputs(6697)) xor (layer0_outputs(9269)));
    layer1_outputs(7279) <= (layer0_outputs(1253)) xor (layer0_outputs(2248));
    layer1_outputs(7280) <= not(layer0_outputs(7686));
    layer1_outputs(7281) <= not((layer0_outputs(8686)) or (layer0_outputs(3082)));
    layer1_outputs(7282) <= not(layer0_outputs(9970)) or (layer0_outputs(6739));
    layer1_outputs(7283) <= layer0_outputs(6207);
    layer1_outputs(7284) <= not((layer0_outputs(7445)) or (layer0_outputs(9460)));
    layer1_outputs(7285) <= not(layer0_outputs(4805));
    layer1_outputs(7286) <= not((layer0_outputs(3364)) and (layer0_outputs(9026)));
    layer1_outputs(7287) <= (layer0_outputs(4155)) and not (layer0_outputs(7296));
    layer1_outputs(7288) <= (layer0_outputs(4673)) xor (layer0_outputs(5788));
    layer1_outputs(7289) <= not((layer0_outputs(4929)) xor (layer0_outputs(2107)));
    layer1_outputs(7290) <= not((layer0_outputs(1889)) and (layer0_outputs(14)));
    layer1_outputs(7291) <= layer0_outputs(6938);
    layer1_outputs(7292) <= not((layer0_outputs(6541)) xor (layer0_outputs(2515)));
    layer1_outputs(7293) <= not(layer0_outputs(5395));
    layer1_outputs(7294) <= (layer0_outputs(3661)) and not (layer0_outputs(100));
    layer1_outputs(7295) <= not((layer0_outputs(132)) or (layer0_outputs(9144)));
    layer1_outputs(7296) <= layer0_outputs(2332);
    layer1_outputs(7297) <= layer0_outputs(8196);
    layer1_outputs(7298) <= not(layer0_outputs(1729)) or (layer0_outputs(4362));
    layer1_outputs(7299) <= layer0_outputs(765);
    layer1_outputs(7300) <= layer0_outputs(5388);
    layer1_outputs(7301) <= not((layer0_outputs(8112)) or (layer0_outputs(2686)));
    layer1_outputs(7302) <= (layer0_outputs(1855)) xor (layer0_outputs(5575));
    layer1_outputs(7303) <= (layer0_outputs(4427)) and not (layer0_outputs(1447));
    layer1_outputs(7304) <= (layer0_outputs(7428)) and (layer0_outputs(14));
    layer1_outputs(7305) <= layer0_outputs(2217);
    layer1_outputs(7306) <= not(layer0_outputs(7177));
    layer1_outputs(7307) <= layer0_outputs(6379);
    layer1_outputs(7308) <= (layer0_outputs(5628)) and not (layer0_outputs(6596));
    layer1_outputs(7309) <= layer0_outputs(3249);
    layer1_outputs(7310) <= not((layer0_outputs(4019)) and (layer0_outputs(9958)));
    layer1_outputs(7311) <= not(layer0_outputs(10224));
    layer1_outputs(7312) <= layer0_outputs(4892);
    layer1_outputs(7313) <= '0';
    layer1_outputs(7314) <= layer0_outputs(6275);
    layer1_outputs(7315) <= not(layer0_outputs(7279));
    layer1_outputs(7316) <= not((layer0_outputs(4445)) or (layer0_outputs(7114)));
    layer1_outputs(7317) <= layer0_outputs(5380);
    layer1_outputs(7318) <= not((layer0_outputs(5114)) xor (layer0_outputs(2851)));
    layer1_outputs(7319) <= not(layer0_outputs(155));
    layer1_outputs(7320) <= (layer0_outputs(8479)) and not (layer0_outputs(3955));
    layer1_outputs(7321) <= (layer0_outputs(5883)) xor (layer0_outputs(9056));
    layer1_outputs(7322) <= (layer0_outputs(6382)) or (layer0_outputs(10195));
    layer1_outputs(7323) <= (layer0_outputs(2803)) and not (layer0_outputs(1524));
    layer1_outputs(7324) <= not(layer0_outputs(5989));
    layer1_outputs(7325) <= not(layer0_outputs(4209));
    layer1_outputs(7326) <= (layer0_outputs(9382)) and not (layer0_outputs(8667));
    layer1_outputs(7327) <= not(layer0_outputs(6574));
    layer1_outputs(7328) <= not(layer0_outputs(4616)) or (layer0_outputs(7929));
    layer1_outputs(7329) <= not(layer0_outputs(3767));
    layer1_outputs(7330) <= not(layer0_outputs(1012));
    layer1_outputs(7331) <= not((layer0_outputs(10023)) xor (layer0_outputs(9777)));
    layer1_outputs(7332) <= not((layer0_outputs(2033)) xor (layer0_outputs(8293)));
    layer1_outputs(7333) <= (layer0_outputs(6062)) and not (layer0_outputs(2554));
    layer1_outputs(7334) <= layer0_outputs(10201);
    layer1_outputs(7335) <= layer0_outputs(7043);
    layer1_outputs(7336) <= layer0_outputs(701);
    layer1_outputs(7337) <= (layer0_outputs(2726)) and not (layer0_outputs(5710));
    layer1_outputs(7338) <= (layer0_outputs(9251)) xor (layer0_outputs(1550));
    layer1_outputs(7339) <= not((layer0_outputs(3116)) and (layer0_outputs(7131)));
    layer1_outputs(7340) <= not((layer0_outputs(7021)) xor (layer0_outputs(2121)));
    layer1_outputs(7341) <= (layer0_outputs(54)) and not (layer0_outputs(9590));
    layer1_outputs(7342) <= '0';
    layer1_outputs(7343) <= layer0_outputs(1471);
    layer1_outputs(7344) <= not((layer0_outputs(8411)) xor (layer0_outputs(1786)));
    layer1_outputs(7345) <= not(layer0_outputs(6397));
    layer1_outputs(7346) <= not(layer0_outputs(4692)) or (layer0_outputs(4234));
    layer1_outputs(7347) <= layer0_outputs(1829);
    layer1_outputs(7348) <= not(layer0_outputs(5239));
    layer1_outputs(7349) <= (layer0_outputs(4587)) and (layer0_outputs(9975));
    layer1_outputs(7350) <= not(layer0_outputs(2270));
    layer1_outputs(7351) <= (layer0_outputs(1619)) and (layer0_outputs(836));
    layer1_outputs(7352) <= (layer0_outputs(7924)) and (layer0_outputs(3929));
    layer1_outputs(7353) <= not((layer0_outputs(2643)) xor (layer0_outputs(2318)));
    layer1_outputs(7354) <= not((layer0_outputs(4902)) xor (layer0_outputs(4243)));
    layer1_outputs(7355) <= '0';
    layer1_outputs(7356) <= layer0_outputs(1256);
    layer1_outputs(7357) <= not((layer0_outputs(8508)) xor (layer0_outputs(9150)));
    layer1_outputs(7358) <= not(layer0_outputs(4389));
    layer1_outputs(7359) <= '0';
    layer1_outputs(7360) <= not((layer0_outputs(4167)) and (layer0_outputs(5864)));
    layer1_outputs(7361) <= '1';
    layer1_outputs(7362) <= not((layer0_outputs(231)) or (layer0_outputs(1945)));
    layer1_outputs(7363) <= not((layer0_outputs(9344)) or (layer0_outputs(6224)));
    layer1_outputs(7364) <= (layer0_outputs(3728)) or (layer0_outputs(3620));
    layer1_outputs(7365) <= (layer0_outputs(1342)) and not (layer0_outputs(8076));
    layer1_outputs(7366) <= layer0_outputs(3249);
    layer1_outputs(7367) <= (layer0_outputs(6613)) or (layer0_outputs(9604));
    layer1_outputs(7368) <= not((layer0_outputs(4315)) and (layer0_outputs(4635)));
    layer1_outputs(7369) <= (layer0_outputs(7680)) and (layer0_outputs(9632));
    layer1_outputs(7370) <= not(layer0_outputs(8365)) or (layer0_outputs(3792));
    layer1_outputs(7371) <= (layer0_outputs(8519)) xor (layer0_outputs(4398));
    layer1_outputs(7372) <= not(layer0_outputs(1699));
    layer1_outputs(7373) <= (layer0_outputs(8395)) and not (layer0_outputs(4992));
    layer1_outputs(7374) <= (layer0_outputs(9790)) and not (layer0_outputs(435));
    layer1_outputs(7375) <= not(layer0_outputs(3440));
    layer1_outputs(7376) <= (layer0_outputs(1284)) or (layer0_outputs(7693));
    layer1_outputs(7377) <= not((layer0_outputs(5195)) xor (layer0_outputs(4017)));
    layer1_outputs(7378) <= layer0_outputs(9748);
    layer1_outputs(7379) <= not((layer0_outputs(7610)) xor (layer0_outputs(3576)));
    layer1_outputs(7380) <= not(layer0_outputs(3861)) or (layer0_outputs(2180));
    layer1_outputs(7381) <= layer0_outputs(8368);
    layer1_outputs(7382) <= not(layer0_outputs(255)) or (layer0_outputs(2473));
    layer1_outputs(7383) <= not(layer0_outputs(158));
    layer1_outputs(7384) <= not(layer0_outputs(4191)) or (layer0_outputs(5590));
    layer1_outputs(7385) <= layer0_outputs(6232);
    layer1_outputs(7386) <= layer0_outputs(8355);
    layer1_outputs(7387) <= (layer0_outputs(3356)) and not (layer0_outputs(3532));
    layer1_outputs(7388) <= not(layer0_outputs(4998));
    layer1_outputs(7389) <= '1';
    layer1_outputs(7390) <= (layer0_outputs(4923)) and not (layer0_outputs(6833));
    layer1_outputs(7391) <= (layer0_outputs(2027)) xor (layer0_outputs(8768));
    layer1_outputs(7392) <= layer0_outputs(4976);
    layer1_outputs(7393) <= layer0_outputs(3323);
    layer1_outputs(7394) <= not(layer0_outputs(5039)) or (layer0_outputs(1108));
    layer1_outputs(7395) <= layer0_outputs(6341);
    layer1_outputs(7396) <= not((layer0_outputs(2466)) and (layer0_outputs(1409)));
    layer1_outputs(7397) <= not(layer0_outputs(5227));
    layer1_outputs(7398) <= not((layer0_outputs(547)) xor (layer0_outputs(1040)));
    layer1_outputs(7399) <= not(layer0_outputs(8688));
    layer1_outputs(7400) <= layer0_outputs(7002);
    layer1_outputs(7401) <= (layer0_outputs(3337)) xor (layer0_outputs(4930));
    layer1_outputs(7402) <= not((layer0_outputs(1279)) and (layer0_outputs(6198)));
    layer1_outputs(7403) <= not(layer0_outputs(1761));
    layer1_outputs(7404) <= not(layer0_outputs(6664));
    layer1_outputs(7405) <= (layer0_outputs(9889)) xor (layer0_outputs(3720));
    layer1_outputs(7406) <= (layer0_outputs(8428)) and not (layer0_outputs(9347));
    layer1_outputs(7407) <= not(layer0_outputs(5912)) or (layer0_outputs(6840));
    layer1_outputs(7408) <= layer0_outputs(2221);
    layer1_outputs(7409) <= not((layer0_outputs(4869)) xor (layer0_outputs(8791)));
    layer1_outputs(7410) <= layer0_outputs(6177);
    layer1_outputs(7411) <= (layer0_outputs(6264)) and (layer0_outputs(2498));
    layer1_outputs(7412) <= (layer0_outputs(7400)) xor (layer0_outputs(664));
    layer1_outputs(7413) <= not(layer0_outputs(6149)) or (layer0_outputs(8058));
    layer1_outputs(7414) <= not(layer0_outputs(3468));
    layer1_outputs(7415) <= layer0_outputs(5953);
    layer1_outputs(7416) <= not((layer0_outputs(4132)) xor (layer0_outputs(3132)));
    layer1_outputs(7417) <= (layer0_outputs(9209)) and not (layer0_outputs(6009));
    layer1_outputs(7418) <= not(layer0_outputs(6342));
    layer1_outputs(7419) <= layer0_outputs(6987);
    layer1_outputs(7420) <= not(layer0_outputs(5899)) or (layer0_outputs(6315));
    layer1_outputs(7421) <= layer0_outputs(7908);
    layer1_outputs(7422) <= layer0_outputs(6119);
    layer1_outputs(7423) <= layer0_outputs(9432);
    layer1_outputs(7424) <= not((layer0_outputs(680)) and (layer0_outputs(8950)));
    layer1_outputs(7425) <= not(layer0_outputs(3208));
    layer1_outputs(7426) <= not((layer0_outputs(2145)) xor (layer0_outputs(8588)));
    layer1_outputs(7427) <= not((layer0_outputs(3820)) or (layer0_outputs(3463)));
    layer1_outputs(7428) <= not((layer0_outputs(7094)) xor (layer0_outputs(4062)));
    layer1_outputs(7429) <= not(layer0_outputs(9949));
    layer1_outputs(7430) <= layer0_outputs(8969);
    layer1_outputs(7431) <= layer0_outputs(5158);
    layer1_outputs(7432) <= not(layer0_outputs(3215)) or (layer0_outputs(968));
    layer1_outputs(7433) <= not((layer0_outputs(4141)) and (layer0_outputs(6392)));
    layer1_outputs(7434) <= (layer0_outputs(4419)) and (layer0_outputs(9228));
    layer1_outputs(7435) <= not((layer0_outputs(9157)) and (layer0_outputs(7187)));
    layer1_outputs(7436) <= not(layer0_outputs(6824));
    layer1_outputs(7437) <= not(layer0_outputs(2393));
    layer1_outputs(7438) <= layer0_outputs(7178);
    layer1_outputs(7439) <= not(layer0_outputs(6598));
    layer1_outputs(7440) <= not((layer0_outputs(7656)) xor (layer0_outputs(1839)));
    layer1_outputs(7441) <= (layer0_outputs(6402)) or (layer0_outputs(4733));
    layer1_outputs(7442) <= layer0_outputs(2751);
    layer1_outputs(7443) <= not(layer0_outputs(26));
    layer1_outputs(7444) <= not((layer0_outputs(1317)) and (layer0_outputs(226)));
    layer1_outputs(7445) <= not(layer0_outputs(7633));
    layer1_outputs(7446) <= not(layer0_outputs(1681));
    layer1_outputs(7447) <= not((layer0_outputs(4198)) xor (layer0_outputs(5796)));
    layer1_outputs(7448) <= (layer0_outputs(2536)) and not (layer0_outputs(221));
    layer1_outputs(7449) <= not(layer0_outputs(6959)) or (layer0_outputs(1785));
    layer1_outputs(7450) <= layer0_outputs(9902);
    layer1_outputs(7451) <= layer0_outputs(3034);
    layer1_outputs(7452) <= not((layer0_outputs(7463)) and (layer0_outputs(1)));
    layer1_outputs(7453) <= (layer0_outputs(9218)) and not (layer0_outputs(7938));
    layer1_outputs(7454) <= layer0_outputs(9782);
    layer1_outputs(7455) <= not(layer0_outputs(4226)) or (layer0_outputs(10063));
    layer1_outputs(7456) <= (layer0_outputs(4924)) xor (layer0_outputs(3072));
    layer1_outputs(7457) <= (layer0_outputs(6526)) and (layer0_outputs(4516));
    layer1_outputs(7458) <= not(layer0_outputs(7159)) or (layer0_outputs(3686));
    layer1_outputs(7459) <= '1';
    layer1_outputs(7460) <= not((layer0_outputs(2800)) or (layer0_outputs(6544)));
    layer1_outputs(7461) <= (layer0_outputs(1082)) and (layer0_outputs(2684));
    layer1_outputs(7462) <= layer0_outputs(9168);
    layer1_outputs(7463) <= not(layer0_outputs(8621)) or (layer0_outputs(6611));
    layer1_outputs(7464) <= (layer0_outputs(9628)) and (layer0_outputs(7837));
    layer1_outputs(7465) <= (layer0_outputs(670)) and not (layer0_outputs(9073));
    layer1_outputs(7466) <= not((layer0_outputs(3079)) xor (layer0_outputs(4074)));
    layer1_outputs(7467) <= (layer0_outputs(8931)) xor (layer0_outputs(2777));
    layer1_outputs(7468) <= (layer0_outputs(6096)) or (layer0_outputs(8298));
    layer1_outputs(7469) <= not(layer0_outputs(7681));
    layer1_outputs(7470) <= (layer0_outputs(3551)) and not (layer0_outputs(3867));
    layer1_outputs(7471) <= not((layer0_outputs(1702)) xor (layer0_outputs(1153)));
    layer1_outputs(7472) <= layer0_outputs(3945);
    layer1_outputs(7473) <= not(layer0_outputs(7646));
    layer1_outputs(7474) <= (layer0_outputs(9516)) or (layer0_outputs(4034));
    layer1_outputs(7475) <= (layer0_outputs(594)) xor (layer0_outputs(498));
    layer1_outputs(7476) <= not(layer0_outputs(5024));
    layer1_outputs(7477) <= (layer0_outputs(2022)) and not (layer0_outputs(903));
    layer1_outputs(7478) <= not(layer0_outputs(1260));
    layer1_outputs(7479) <= layer0_outputs(1546);
    layer1_outputs(7480) <= not((layer0_outputs(5309)) or (layer0_outputs(7826)));
    layer1_outputs(7481) <= layer0_outputs(6155);
    layer1_outputs(7482) <= layer0_outputs(4063);
    layer1_outputs(7483) <= (layer0_outputs(4276)) and (layer0_outputs(6040));
    layer1_outputs(7484) <= not(layer0_outputs(4542)) or (layer0_outputs(10032));
    layer1_outputs(7485) <= (layer0_outputs(8662)) and (layer0_outputs(8787));
    layer1_outputs(7486) <= not(layer0_outputs(7538));
    layer1_outputs(7487) <= (layer0_outputs(1047)) and not (layer0_outputs(5240));
    layer1_outputs(7488) <= not(layer0_outputs(6291));
    layer1_outputs(7489) <= (layer0_outputs(6005)) and not (layer0_outputs(8671));
    layer1_outputs(7490) <= not(layer0_outputs(5817)) or (layer0_outputs(4371));
    layer1_outputs(7491) <= (layer0_outputs(6761)) or (layer0_outputs(5293));
    layer1_outputs(7492) <= not(layer0_outputs(10235));
    layer1_outputs(7493) <= not(layer0_outputs(3841));
    layer1_outputs(7494) <= not(layer0_outputs(2848));
    layer1_outputs(7495) <= not(layer0_outputs(3578)) or (layer0_outputs(6382));
    layer1_outputs(7496) <= not(layer0_outputs(6655));
    layer1_outputs(7497) <= layer0_outputs(8394);
    layer1_outputs(7498) <= not(layer0_outputs(1309));
    layer1_outputs(7499) <= not(layer0_outputs(9639)) or (layer0_outputs(92));
    layer1_outputs(7500) <= (layer0_outputs(1944)) and not (layer0_outputs(10073));
    layer1_outputs(7501) <= layer0_outputs(3282);
    layer1_outputs(7502) <= not(layer0_outputs(2331));
    layer1_outputs(7503) <= (layer0_outputs(1483)) and not (layer0_outputs(1103));
    layer1_outputs(7504) <= (layer0_outputs(7739)) and (layer0_outputs(2310));
    layer1_outputs(7505) <= (layer0_outputs(966)) xor (layer0_outputs(1248));
    layer1_outputs(7506) <= not(layer0_outputs(1885)) or (layer0_outputs(8678));
    layer1_outputs(7507) <= (layer0_outputs(1025)) xor (layer0_outputs(2142));
    layer1_outputs(7508) <= not(layer0_outputs(5228)) or (layer0_outputs(2864));
    layer1_outputs(7509) <= (layer0_outputs(426)) xor (layer0_outputs(4384));
    layer1_outputs(7510) <= not((layer0_outputs(8823)) or (layer0_outputs(2106)));
    layer1_outputs(7511) <= not(layer0_outputs(9904));
    layer1_outputs(7512) <= layer0_outputs(5508);
    layer1_outputs(7513) <= layer0_outputs(5133);
    layer1_outputs(7514) <= layer0_outputs(9601);
    layer1_outputs(7515) <= not((layer0_outputs(8780)) xor (layer0_outputs(7982)));
    layer1_outputs(7516) <= layer0_outputs(5225);
    layer1_outputs(7517) <= layer0_outputs(9849);
    layer1_outputs(7518) <= '1';
    layer1_outputs(7519) <= not(layer0_outputs(7274));
    layer1_outputs(7520) <= not((layer0_outputs(9591)) or (layer0_outputs(5869)));
    layer1_outputs(7521) <= layer0_outputs(2572);
    layer1_outputs(7522) <= layer0_outputs(955);
    layer1_outputs(7523) <= not(layer0_outputs(9170)) or (layer0_outputs(6565));
    layer1_outputs(7524) <= (layer0_outputs(1902)) and not (layer0_outputs(7296));
    layer1_outputs(7525) <= not(layer0_outputs(1710)) or (layer0_outputs(905));
    layer1_outputs(7526) <= (layer0_outputs(9601)) and not (layer0_outputs(4287));
    layer1_outputs(7527) <= not(layer0_outputs(9156));
    layer1_outputs(7528) <= not((layer0_outputs(9017)) xor (layer0_outputs(2688)));
    layer1_outputs(7529) <= not(layer0_outputs(8501)) or (layer0_outputs(4800));
    layer1_outputs(7530) <= not((layer0_outputs(5480)) and (layer0_outputs(9095)));
    layer1_outputs(7531) <= not(layer0_outputs(5917)) or (layer0_outputs(2624));
    layer1_outputs(7532) <= layer0_outputs(1462);
    layer1_outputs(7533) <= (layer0_outputs(7524)) and not (layer0_outputs(3466));
    layer1_outputs(7534) <= layer0_outputs(4648);
    layer1_outputs(7535) <= not((layer0_outputs(6996)) and (layer0_outputs(8618)));
    layer1_outputs(7536) <= (layer0_outputs(6566)) xor (layer0_outputs(9110));
    layer1_outputs(7537) <= not(layer0_outputs(472)) or (layer0_outputs(9361));
    layer1_outputs(7538) <= not((layer0_outputs(2252)) xor (layer0_outputs(5662)));
    layer1_outputs(7539) <= not(layer0_outputs(1570));
    layer1_outputs(7540) <= (layer0_outputs(2029)) and (layer0_outputs(2063));
    layer1_outputs(7541) <= not(layer0_outputs(3684));
    layer1_outputs(7542) <= (layer0_outputs(1455)) and not (layer0_outputs(1559));
    layer1_outputs(7543) <= not((layer0_outputs(6101)) xor (layer0_outputs(1481)));
    layer1_outputs(7544) <= layer0_outputs(10153);
    layer1_outputs(7545) <= (layer0_outputs(3284)) and not (layer0_outputs(499));
    layer1_outputs(7546) <= not(layer0_outputs(9121));
    layer1_outputs(7547) <= not(layer0_outputs(8415));
    layer1_outputs(7548) <= not(layer0_outputs(8875));
    layer1_outputs(7549) <= not(layer0_outputs(294));
    layer1_outputs(7550) <= '0';
    layer1_outputs(7551) <= not(layer0_outputs(7434)) or (layer0_outputs(2911));
    layer1_outputs(7552) <= not((layer0_outputs(4364)) xor (layer0_outputs(2778)));
    layer1_outputs(7553) <= layer0_outputs(3834);
    layer1_outputs(7554) <= layer0_outputs(4353);
    layer1_outputs(7555) <= (layer0_outputs(8061)) xor (layer0_outputs(2161));
    layer1_outputs(7556) <= (layer0_outputs(3965)) and (layer0_outputs(3430));
    layer1_outputs(7557) <= (layer0_outputs(212)) and (layer0_outputs(1490));
    layer1_outputs(7558) <= '0';
    layer1_outputs(7559) <= layer0_outputs(8535);
    layer1_outputs(7560) <= not(layer0_outputs(8210)) or (layer0_outputs(6531));
    layer1_outputs(7561) <= layer0_outputs(1358);
    layer1_outputs(7562) <= (layer0_outputs(5258)) and not (layer0_outputs(257));
    layer1_outputs(7563) <= not(layer0_outputs(1238));
    layer1_outputs(7564) <= not(layer0_outputs(6932));
    layer1_outputs(7565) <= layer0_outputs(376);
    layer1_outputs(7566) <= (layer0_outputs(2338)) or (layer0_outputs(7198));
    layer1_outputs(7567) <= not(layer0_outputs(5948));
    layer1_outputs(7568) <= (layer0_outputs(2464)) and not (layer0_outputs(1988));
    layer1_outputs(7569) <= '1';
    layer1_outputs(7570) <= not((layer0_outputs(3019)) and (layer0_outputs(10016)));
    layer1_outputs(7571) <= not(layer0_outputs(3458));
    layer1_outputs(7572) <= not((layer0_outputs(3107)) xor (layer0_outputs(8750)));
    layer1_outputs(7573) <= layer0_outputs(5754);
    layer1_outputs(7574) <= layer0_outputs(4464);
    layer1_outputs(7575) <= (layer0_outputs(8654)) or (layer0_outputs(3265));
    layer1_outputs(7576) <= not((layer0_outputs(2926)) or (layer0_outputs(5555)));
    layer1_outputs(7577) <= not((layer0_outputs(5573)) xor (layer0_outputs(5845)));
    layer1_outputs(7578) <= (layer0_outputs(5142)) or (layer0_outputs(8407));
    layer1_outputs(7579) <= layer0_outputs(5276);
    layer1_outputs(7580) <= (layer0_outputs(6609)) and not (layer0_outputs(7932));
    layer1_outputs(7581) <= layer0_outputs(5202);
    layer1_outputs(7582) <= not((layer0_outputs(8035)) or (layer0_outputs(5089)));
    layer1_outputs(7583) <= not((layer0_outputs(1713)) or (layer0_outputs(4725)));
    layer1_outputs(7584) <= not(layer0_outputs(4218));
    layer1_outputs(7585) <= not(layer0_outputs(10130));
    layer1_outputs(7586) <= (layer0_outputs(2031)) and not (layer0_outputs(7863));
    layer1_outputs(7587) <= not((layer0_outputs(4662)) and (layer0_outputs(9355)));
    layer1_outputs(7588) <= layer0_outputs(5973);
    layer1_outputs(7589) <= not(layer0_outputs(4926));
    layer1_outputs(7590) <= not((layer0_outputs(8698)) and (layer0_outputs(4434)));
    layer1_outputs(7591) <= layer0_outputs(5286);
    layer1_outputs(7592) <= not(layer0_outputs(2635)) or (layer0_outputs(8263));
    layer1_outputs(7593) <= (layer0_outputs(5364)) and (layer0_outputs(2768));
    layer1_outputs(7594) <= not(layer0_outputs(3702));
    layer1_outputs(7595) <= (layer0_outputs(1415)) and (layer0_outputs(2818));
    layer1_outputs(7596) <= (layer0_outputs(6150)) and not (layer0_outputs(8708));
    layer1_outputs(7597) <= (layer0_outputs(8417)) or (layer0_outputs(571));
    layer1_outputs(7598) <= not(layer0_outputs(9694));
    layer1_outputs(7599) <= '0';
    layer1_outputs(7600) <= layer0_outputs(939);
    layer1_outputs(7601) <= (layer0_outputs(9788)) and (layer0_outputs(5984));
    layer1_outputs(7602) <= layer0_outputs(9849);
    layer1_outputs(7603) <= not(layer0_outputs(5833));
    layer1_outputs(7604) <= layer0_outputs(286);
    layer1_outputs(7605) <= not((layer0_outputs(52)) or (layer0_outputs(545)));
    layer1_outputs(7606) <= '1';
    layer1_outputs(7607) <= not((layer0_outputs(2716)) and (layer0_outputs(7569)));
    layer1_outputs(7608) <= (layer0_outputs(1706)) and not (layer0_outputs(4993));
    layer1_outputs(7609) <= layer0_outputs(1659);
    layer1_outputs(7610) <= layer0_outputs(7615);
    layer1_outputs(7611) <= (layer0_outputs(9461)) and not (layer0_outputs(4877));
    layer1_outputs(7612) <= (layer0_outputs(9987)) and not (layer0_outputs(1237));
    layer1_outputs(7613) <= not((layer0_outputs(8539)) and (layer0_outputs(8743)));
    layer1_outputs(7614) <= (layer0_outputs(7121)) or (layer0_outputs(3078));
    layer1_outputs(7615) <= not(layer0_outputs(4927));
    layer1_outputs(7616) <= not(layer0_outputs(9309)) or (layer0_outputs(9243));
    layer1_outputs(7617) <= '1';
    layer1_outputs(7618) <= layer0_outputs(127);
    layer1_outputs(7619) <= layer0_outputs(9310);
    layer1_outputs(7620) <= layer0_outputs(10145);
    layer1_outputs(7621) <= (layer0_outputs(3650)) and not (layer0_outputs(3639));
    layer1_outputs(7622) <= not((layer0_outputs(6272)) or (layer0_outputs(614)));
    layer1_outputs(7623) <= not((layer0_outputs(7403)) and (layer0_outputs(8242)));
    layer1_outputs(7624) <= not(layer0_outputs(6078));
    layer1_outputs(7625) <= (layer0_outputs(6683)) and not (layer0_outputs(4288));
    layer1_outputs(7626) <= (layer0_outputs(2789)) and not (layer0_outputs(6266));
    layer1_outputs(7627) <= (layer0_outputs(4966)) or (layer0_outputs(2622));
    layer1_outputs(7628) <= layer0_outputs(9440);
    layer1_outputs(7629) <= layer0_outputs(5427);
    layer1_outputs(7630) <= not(layer0_outputs(6023));
    layer1_outputs(7631) <= (layer0_outputs(6232)) or (layer0_outputs(2357));
    layer1_outputs(7632) <= '1';
    layer1_outputs(7633) <= not(layer0_outputs(9162));
    layer1_outputs(7634) <= not(layer0_outputs(5674));
    layer1_outputs(7635) <= not(layer0_outputs(2141)) or (layer0_outputs(1576));
    layer1_outputs(7636) <= layer0_outputs(4238);
    layer1_outputs(7637) <= layer0_outputs(8046);
    layer1_outputs(7638) <= (layer0_outputs(7045)) or (layer0_outputs(4076));
    layer1_outputs(7639) <= (layer0_outputs(6830)) and (layer0_outputs(4788));
    layer1_outputs(7640) <= not((layer0_outputs(9262)) xor (layer0_outputs(2774)));
    layer1_outputs(7641) <= not(layer0_outputs(7877));
    layer1_outputs(7642) <= not(layer0_outputs(4533));
    layer1_outputs(7643) <= not(layer0_outputs(1554)) or (layer0_outputs(2360));
    layer1_outputs(7644) <= layer0_outputs(1469);
    layer1_outputs(7645) <= not(layer0_outputs(207));
    layer1_outputs(7646) <= not(layer0_outputs(9900)) or (layer0_outputs(5580));
    layer1_outputs(7647) <= not(layer0_outputs(117)) or (layer0_outputs(7516));
    layer1_outputs(7648) <= (layer0_outputs(7809)) xor (layer0_outputs(10028));
    layer1_outputs(7649) <= (layer0_outputs(1673)) and not (layer0_outputs(7564));
    layer1_outputs(7650) <= not((layer0_outputs(216)) or (layer0_outputs(8019)));
    layer1_outputs(7651) <= (layer0_outputs(848)) and not (layer0_outputs(6942));
    layer1_outputs(7652) <= '1';
    layer1_outputs(7653) <= (layer0_outputs(7484)) and not (layer0_outputs(3762));
    layer1_outputs(7654) <= layer0_outputs(7239);
    layer1_outputs(7655) <= (layer0_outputs(1159)) xor (layer0_outputs(9131));
    layer1_outputs(7656) <= not(layer0_outputs(4175));
    layer1_outputs(7657) <= not((layer0_outputs(7651)) and (layer0_outputs(6865)));
    layer1_outputs(7658) <= (layer0_outputs(4175)) xor (layer0_outputs(4705));
    layer1_outputs(7659) <= (layer0_outputs(1167)) and (layer0_outputs(3118));
    layer1_outputs(7660) <= layer0_outputs(2355);
    layer1_outputs(7661) <= not(layer0_outputs(5879)) or (layer0_outputs(6463));
    layer1_outputs(7662) <= not((layer0_outputs(2489)) or (layer0_outputs(9440)));
    layer1_outputs(7663) <= (layer0_outputs(9731)) xor (layer0_outputs(2121));
    layer1_outputs(7664) <= layer0_outputs(7468);
    layer1_outputs(7665) <= not(layer0_outputs(9395));
    layer1_outputs(7666) <= not(layer0_outputs(1650));
    layer1_outputs(7667) <= not(layer0_outputs(2238));
    layer1_outputs(7668) <= (layer0_outputs(4502)) or (layer0_outputs(8393));
    layer1_outputs(7669) <= '0';
    layer1_outputs(7670) <= (layer0_outputs(3058)) xor (layer0_outputs(7308));
    layer1_outputs(7671) <= not((layer0_outputs(4604)) or (layer0_outputs(8040)));
    layer1_outputs(7672) <= not((layer0_outputs(1933)) xor (layer0_outputs(1598)));
    layer1_outputs(7673) <= not((layer0_outputs(6086)) and (layer0_outputs(4619)));
    layer1_outputs(7674) <= not(layer0_outputs(9939)) or (layer0_outputs(7325));
    layer1_outputs(7675) <= not(layer0_outputs(4503));
    layer1_outputs(7676) <= (layer0_outputs(1535)) and not (layer0_outputs(1798));
    layer1_outputs(7677) <= layer0_outputs(9722);
    layer1_outputs(7678) <= not(layer0_outputs(3473));
    layer1_outputs(7679) <= layer0_outputs(1420);
    layer1_outputs(7680) <= (layer0_outputs(2438)) and (layer0_outputs(1777));
    layer1_outputs(7681) <= layer0_outputs(6737);
    layer1_outputs(7682) <= (layer0_outputs(7362)) and not (layer0_outputs(5485));
    layer1_outputs(7683) <= not(layer0_outputs(3644));
    layer1_outputs(7684) <= not(layer0_outputs(15));
    layer1_outputs(7685) <= layer0_outputs(9925);
    layer1_outputs(7686) <= not(layer0_outputs(3997));
    layer1_outputs(7687) <= layer0_outputs(8721);
    layer1_outputs(7688) <= layer0_outputs(5782);
    layer1_outputs(7689) <= not(layer0_outputs(691));
    layer1_outputs(7690) <= (layer0_outputs(774)) and not (layer0_outputs(4934));
    layer1_outputs(7691) <= (layer0_outputs(7525)) xor (layer0_outputs(9348));
    layer1_outputs(7692) <= not((layer0_outputs(8830)) xor (layer0_outputs(7653)));
    layer1_outputs(7693) <= (layer0_outputs(10060)) and not (layer0_outputs(6700));
    layer1_outputs(7694) <= not((layer0_outputs(5569)) and (layer0_outputs(1081)));
    layer1_outputs(7695) <= layer0_outputs(384);
    layer1_outputs(7696) <= not((layer0_outputs(417)) and (layer0_outputs(3509)));
    layer1_outputs(7697) <= not(layer0_outputs(4828)) or (layer0_outputs(140));
    layer1_outputs(7698) <= (layer0_outputs(7012)) xor (layer0_outputs(7417));
    layer1_outputs(7699) <= (layer0_outputs(2039)) and not (layer0_outputs(7549));
    layer1_outputs(7700) <= (layer0_outputs(8324)) and (layer0_outputs(8658));
    layer1_outputs(7701) <= not((layer0_outputs(3066)) xor (layer0_outputs(8352)));
    layer1_outputs(7702) <= not(layer0_outputs(5462)) or (layer0_outputs(4433));
    layer1_outputs(7703) <= layer0_outputs(6014);
    layer1_outputs(7704) <= not((layer0_outputs(9511)) and (layer0_outputs(8571)));
    layer1_outputs(7705) <= not(layer0_outputs(7453));
    layer1_outputs(7706) <= not(layer0_outputs(9313));
    layer1_outputs(7707) <= layer0_outputs(6281);
    layer1_outputs(7708) <= layer0_outputs(2777);
    layer1_outputs(7709) <= not((layer0_outputs(7825)) or (layer0_outputs(3587)));
    layer1_outputs(7710) <= layer0_outputs(5349);
    layer1_outputs(7711) <= not((layer0_outputs(7614)) and (layer0_outputs(3311)));
    layer1_outputs(7712) <= layer0_outputs(7406);
    layer1_outputs(7713) <= (layer0_outputs(4743)) and (layer0_outputs(5257));
    layer1_outputs(7714) <= not((layer0_outputs(8945)) and (layer0_outputs(9022)));
    layer1_outputs(7715) <= (layer0_outputs(3122)) or (layer0_outputs(8974));
    layer1_outputs(7716) <= (layer0_outputs(7820)) and not (layer0_outputs(710));
    layer1_outputs(7717) <= not((layer0_outputs(3425)) or (layer0_outputs(6183)));
    layer1_outputs(7718) <= not(layer0_outputs(2570));
    layer1_outputs(7719) <= (layer0_outputs(263)) and (layer0_outputs(2288));
    layer1_outputs(7720) <= '0';
    layer1_outputs(7721) <= not((layer0_outputs(111)) or (layer0_outputs(7155)));
    layer1_outputs(7722) <= not(layer0_outputs(2542));
    layer1_outputs(7723) <= (layer0_outputs(1271)) and not (layer0_outputs(3159));
    layer1_outputs(7724) <= not(layer0_outputs(574));
    layer1_outputs(7725) <= layer0_outputs(896);
    layer1_outputs(7726) <= not(layer0_outputs(9117));
    layer1_outputs(7727) <= not(layer0_outputs(6875));
    layer1_outputs(7728) <= not(layer0_outputs(9333));
    layer1_outputs(7729) <= (layer0_outputs(8496)) xor (layer0_outputs(990));
    layer1_outputs(7730) <= (layer0_outputs(4195)) and (layer0_outputs(6777));
    layer1_outputs(7731) <= (layer0_outputs(6429)) and not (layer0_outputs(9658));
    layer1_outputs(7732) <= layer0_outputs(1468);
    layer1_outputs(7733) <= '1';
    layer1_outputs(7734) <= not((layer0_outputs(6762)) xor (layer0_outputs(5803)));
    layer1_outputs(7735) <= not(layer0_outputs(6713)) or (layer0_outputs(3698));
    layer1_outputs(7736) <= layer0_outputs(9815);
    layer1_outputs(7737) <= layer0_outputs(7450);
    layer1_outputs(7738) <= not((layer0_outputs(7608)) and (layer0_outputs(9124)));
    layer1_outputs(7739) <= layer0_outputs(3187);
    layer1_outputs(7740) <= not(layer0_outputs(8785));
    layer1_outputs(7741) <= (layer0_outputs(1096)) and (layer0_outputs(5054));
    layer1_outputs(7742) <= layer0_outputs(7711);
    layer1_outputs(7743) <= not(layer0_outputs(8514));
    layer1_outputs(7744) <= not(layer0_outputs(2459));
    layer1_outputs(7745) <= layer0_outputs(5957);
    layer1_outputs(7746) <= not((layer0_outputs(4555)) xor (layer0_outputs(9371)));
    layer1_outputs(7747) <= (layer0_outputs(4594)) or (layer0_outputs(7579));
    layer1_outputs(7748) <= not(layer0_outputs(3266));
    layer1_outputs(7749) <= layer0_outputs(3590);
    layer1_outputs(7750) <= not((layer0_outputs(7674)) xor (layer0_outputs(1295)));
    layer1_outputs(7751) <= not(layer0_outputs(2653));
    layer1_outputs(7752) <= (layer0_outputs(8531)) and (layer0_outputs(812));
    layer1_outputs(7753) <= layer0_outputs(5884);
    layer1_outputs(7754) <= not((layer0_outputs(427)) and (layer0_outputs(189)));
    layer1_outputs(7755) <= (layer0_outputs(7512)) xor (layer0_outputs(5411));
    layer1_outputs(7756) <= (layer0_outputs(508)) and not (layer0_outputs(6740));
    layer1_outputs(7757) <= not(layer0_outputs(8418)) or (layer0_outputs(2401));
    layer1_outputs(7758) <= not((layer0_outputs(8764)) and (layer0_outputs(5258)));
    layer1_outputs(7759) <= not(layer0_outputs(3517));
    layer1_outputs(7760) <= not(layer0_outputs(3782));
    layer1_outputs(7761) <= layer0_outputs(2927);
    layer1_outputs(7762) <= (layer0_outputs(6038)) and not (layer0_outputs(8464));
    layer1_outputs(7763) <= (layer0_outputs(4782)) and not (layer0_outputs(5682));
    layer1_outputs(7764) <= (layer0_outputs(319)) and (layer0_outputs(6720));
    layer1_outputs(7765) <= not(layer0_outputs(7662)) or (layer0_outputs(1809));
    layer1_outputs(7766) <= '0';
    layer1_outputs(7767) <= not((layer0_outputs(3540)) xor (layer0_outputs(4006)));
    layer1_outputs(7768) <= '1';
    layer1_outputs(7769) <= not(layer0_outputs(7410));
    layer1_outputs(7770) <= not(layer0_outputs(5249)) or (layer0_outputs(7289));
    layer1_outputs(7771) <= not((layer0_outputs(368)) xor (layer0_outputs(8651)));
    layer1_outputs(7772) <= not(layer0_outputs(9892));
    layer1_outputs(7773) <= layer0_outputs(492);
    layer1_outputs(7774) <= not(layer0_outputs(5927)) or (layer0_outputs(8789));
    layer1_outputs(7775) <= not((layer0_outputs(6862)) or (layer0_outputs(6216)));
    layer1_outputs(7776) <= (layer0_outputs(1236)) or (layer0_outputs(5455));
    layer1_outputs(7777) <= not(layer0_outputs(4093));
    layer1_outputs(7778) <= layer0_outputs(1346);
    layer1_outputs(7779) <= (layer0_outputs(5705)) and not (layer0_outputs(842));
    layer1_outputs(7780) <= (layer0_outputs(9041)) and not (layer0_outputs(4915));
    layer1_outputs(7781) <= (layer0_outputs(8012)) and not (layer0_outputs(6779));
    layer1_outputs(7782) <= not(layer0_outputs(8576));
    layer1_outputs(7783) <= not(layer0_outputs(4611));
    layer1_outputs(7784) <= (layer0_outputs(2172)) and not (layer0_outputs(5223));
    layer1_outputs(7785) <= (layer0_outputs(1703)) xor (layer0_outputs(561));
    layer1_outputs(7786) <= not(layer0_outputs(8284)) or (layer0_outputs(1572));
    layer1_outputs(7787) <= (layer0_outputs(1243)) and not (layer0_outputs(10063));
    layer1_outputs(7788) <= layer0_outputs(6118);
    layer1_outputs(7789) <= (layer0_outputs(218)) xor (layer0_outputs(1765));
    layer1_outputs(7790) <= not(layer0_outputs(5307));
    layer1_outputs(7791) <= layer0_outputs(5100);
    layer1_outputs(7792) <= (layer0_outputs(7306)) and not (layer0_outputs(3984));
    layer1_outputs(7793) <= (layer0_outputs(4118)) and not (layer0_outputs(4952));
    layer1_outputs(7794) <= not(layer0_outputs(8849));
    layer1_outputs(7795) <= layer0_outputs(7320);
    layer1_outputs(7796) <= layer0_outputs(6971);
    layer1_outputs(7797) <= (layer0_outputs(2720)) or (layer0_outputs(6503));
    layer1_outputs(7798) <= '0';
    layer1_outputs(7799) <= layer0_outputs(6663);
    layer1_outputs(7800) <= '1';
    layer1_outputs(7801) <= not((layer0_outputs(742)) xor (layer0_outputs(834)));
    layer1_outputs(7802) <= not(layer0_outputs(10040)) or (layer0_outputs(8246));
    layer1_outputs(7803) <= (layer0_outputs(10140)) and (layer0_outputs(5500));
    layer1_outputs(7804) <= not(layer0_outputs(8032));
    layer1_outputs(7805) <= (layer0_outputs(9513)) and not (layer0_outputs(6102));
    layer1_outputs(7806) <= (layer0_outputs(1266)) and (layer0_outputs(8544));
    layer1_outputs(7807) <= layer0_outputs(390);
    layer1_outputs(7808) <= not(layer0_outputs(764));
    layer1_outputs(7809) <= (layer0_outputs(5304)) or (layer0_outputs(6280));
    layer1_outputs(7810) <= (layer0_outputs(4938)) and not (layer0_outputs(8390));
    layer1_outputs(7811) <= (layer0_outputs(9408)) or (layer0_outputs(4827));
    layer1_outputs(7812) <= not(layer0_outputs(4417));
    layer1_outputs(7813) <= '1';
    layer1_outputs(7814) <= (layer0_outputs(6414)) and not (layer0_outputs(9471));
    layer1_outputs(7815) <= not(layer0_outputs(143)) or (layer0_outputs(9972));
    layer1_outputs(7816) <= not(layer0_outputs(3747)) or (layer0_outputs(8457));
    layer1_outputs(7817) <= not(layer0_outputs(4352));
    layer1_outputs(7818) <= (layer0_outputs(2124)) xor (layer0_outputs(6881));
    layer1_outputs(7819) <= not((layer0_outputs(4937)) xor (layer0_outputs(1269)));
    layer1_outputs(7820) <= not(layer0_outputs(2173)) or (layer0_outputs(9227));
    layer1_outputs(7821) <= layer0_outputs(2644);
    layer1_outputs(7822) <= not(layer0_outputs(4955));
    layer1_outputs(7823) <= not((layer0_outputs(7244)) and (layer0_outputs(1123)));
    layer1_outputs(7824) <= (layer0_outputs(5290)) and (layer0_outputs(8610));
    layer1_outputs(7825) <= not(layer0_outputs(4345));
    layer1_outputs(7826) <= layer0_outputs(7485);
    layer1_outputs(7827) <= layer0_outputs(8038);
    layer1_outputs(7828) <= (layer0_outputs(9998)) xor (layer0_outputs(1762));
    layer1_outputs(7829) <= (layer0_outputs(5323)) or (layer0_outputs(1545));
    layer1_outputs(7830) <= not((layer0_outputs(6851)) or (layer0_outputs(4043)));
    layer1_outputs(7831) <= not(layer0_outputs(9580));
    layer1_outputs(7832) <= (layer0_outputs(4093)) and not (layer0_outputs(5018));
    layer1_outputs(7833) <= layer0_outputs(3041);
    layer1_outputs(7834) <= not((layer0_outputs(4190)) and (layer0_outputs(3781)));
    layer1_outputs(7835) <= layer0_outputs(7838);
    layer1_outputs(7836) <= not((layer0_outputs(705)) and (layer0_outputs(683)));
    layer1_outputs(7837) <= not(layer0_outputs(3547));
    layer1_outputs(7838) <= (layer0_outputs(7961)) or (layer0_outputs(3333));
    layer1_outputs(7839) <= not((layer0_outputs(2916)) xor (layer0_outputs(1904)));
    layer1_outputs(7840) <= (layer0_outputs(5681)) xor (layer0_outputs(2976));
    layer1_outputs(7841) <= (layer0_outputs(7780)) or (layer0_outputs(6406));
    layer1_outputs(7842) <= (layer0_outputs(9893)) and not (layer0_outputs(9685));
    layer1_outputs(7843) <= not((layer0_outputs(2854)) and (layer0_outputs(1348)));
    layer1_outputs(7844) <= (layer0_outputs(7640)) xor (layer0_outputs(6606));
    layer1_outputs(7845) <= '0';
    layer1_outputs(7846) <= layer0_outputs(9840);
    layer1_outputs(7847) <= not(layer0_outputs(3653));
    layer1_outputs(7848) <= not(layer0_outputs(3279));
    layer1_outputs(7849) <= layer0_outputs(7805);
    layer1_outputs(7850) <= layer0_outputs(2278);
    layer1_outputs(7851) <= not((layer0_outputs(843)) xor (layer0_outputs(4941)));
    layer1_outputs(7852) <= layer0_outputs(2936);
    layer1_outputs(7853) <= not(layer0_outputs(860));
    layer1_outputs(7854) <= not(layer0_outputs(9894));
    layer1_outputs(7855) <= layer0_outputs(7998);
    layer1_outputs(7856) <= (layer0_outputs(4757)) and not (layer0_outputs(930));
    layer1_outputs(7857) <= not(layer0_outputs(5982)) or (layer0_outputs(8680));
    layer1_outputs(7858) <= (layer0_outputs(2356)) or (layer0_outputs(3587));
    layer1_outputs(7859) <= (layer0_outputs(144)) and not (layer0_outputs(5581));
    layer1_outputs(7860) <= not((layer0_outputs(10163)) or (layer0_outputs(7342)));
    layer1_outputs(7861) <= not(layer0_outputs(5801)) or (layer0_outputs(5129));
    layer1_outputs(7862) <= layer0_outputs(8608);
    layer1_outputs(7863) <= '1';
    layer1_outputs(7864) <= (layer0_outputs(6509)) and not (layer0_outputs(5311));
    layer1_outputs(7865) <= not((layer0_outputs(5388)) or (layer0_outputs(6828)));
    layer1_outputs(7866) <= (layer0_outputs(7572)) and not (layer0_outputs(7290));
    layer1_outputs(7867) <= layer0_outputs(3693);
    layer1_outputs(7868) <= not(layer0_outputs(2887));
    layer1_outputs(7869) <= not(layer0_outputs(758)) or (layer0_outputs(3618));
    layer1_outputs(7870) <= (layer0_outputs(3269)) and (layer0_outputs(1365));
    layer1_outputs(7871) <= not(layer0_outputs(9304));
    layer1_outputs(7872) <= layer0_outputs(4363);
    layer1_outputs(7873) <= (layer0_outputs(2240)) or (layer0_outputs(959));
    layer1_outputs(7874) <= not(layer0_outputs(5994));
    layer1_outputs(7875) <= (layer0_outputs(4419)) xor (layer0_outputs(9380));
    layer1_outputs(7876) <= not(layer0_outputs(9999));
    layer1_outputs(7877) <= not(layer0_outputs(6537)) or (layer0_outputs(370));
    layer1_outputs(7878) <= not(layer0_outputs(722));
    layer1_outputs(7879) <= not(layer0_outputs(4463));
    layer1_outputs(7880) <= not(layer0_outputs(6335)) or (layer0_outputs(6285));
    layer1_outputs(7881) <= not((layer0_outputs(9786)) or (layer0_outputs(6935)));
    layer1_outputs(7882) <= not(layer0_outputs(6871));
    layer1_outputs(7883) <= (layer0_outputs(9222)) xor (layer0_outputs(4956));
    layer1_outputs(7884) <= (layer0_outputs(9442)) or (layer0_outputs(5493));
    layer1_outputs(7885) <= (layer0_outputs(6668)) and (layer0_outputs(4797));
    layer1_outputs(7886) <= (layer0_outputs(7881)) and (layer0_outputs(4220));
    layer1_outputs(7887) <= not(layer0_outputs(1022)) or (layer0_outputs(2619));
    layer1_outputs(7888) <= not((layer0_outputs(5622)) or (layer0_outputs(405)));
    layer1_outputs(7889) <= (layer0_outputs(9718)) xor (layer0_outputs(5424));
    layer1_outputs(7890) <= not(layer0_outputs(1579));
    layer1_outputs(7891) <= layer0_outputs(7101);
    layer1_outputs(7892) <= not((layer0_outputs(3375)) or (layer0_outputs(5823)));
    layer1_outputs(7893) <= layer0_outputs(1097);
    layer1_outputs(7894) <= not(layer0_outputs(621));
    layer1_outputs(7895) <= layer0_outputs(366);
    layer1_outputs(7896) <= not(layer0_outputs(3121)) or (layer0_outputs(1226));
    layer1_outputs(7897) <= (layer0_outputs(8140)) or (layer0_outputs(9230));
    layer1_outputs(7898) <= not(layer0_outputs(4056));
    layer1_outputs(7899) <= not((layer0_outputs(2074)) xor (layer0_outputs(1323)));
    layer1_outputs(7900) <= layer0_outputs(6489);
    layer1_outputs(7901) <= (layer0_outputs(8364)) and not (layer0_outputs(5214));
    layer1_outputs(7902) <= (layer0_outputs(5294)) or (layer0_outputs(6322));
    layer1_outputs(7903) <= (layer0_outputs(3696)) and (layer0_outputs(4149));
    layer1_outputs(7904) <= not((layer0_outputs(2635)) and (layer0_outputs(9922)));
    layer1_outputs(7905) <= (layer0_outputs(814)) and not (layer0_outputs(5245));
    layer1_outputs(7906) <= not(layer0_outputs(5237));
    layer1_outputs(7907) <= layer0_outputs(4595);
    layer1_outputs(7908) <= (layer0_outputs(1571)) or (layer0_outputs(8516));
    layer1_outputs(7909) <= layer0_outputs(102);
    layer1_outputs(7910) <= not((layer0_outputs(9939)) xor (layer0_outputs(2034)));
    layer1_outputs(7911) <= (layer0_outputs(9173)) and (layer0_outputs(557));
    layer1_outputs(7912) <= layer0_outputs(8659);
    layer1_outputs(7913) <= '0';
    layer1_outputs(7914) <= (layer0_outputs(4977)) and not (layer0_outputs(5370));
    layer1_outputs(7915) <= not((layer0_outputs(930)) or (layer0_outputs(5134)));
    layer1_outputs(7916) <= not(layer0_outputs(8649));
    layer1_outputs(7917) <= (layer0_outputs(4176)) xor (layer0_outputs(3877));
    layer1_outputs(7918) <= layer0_outputs(3391);
    layer1_outputs(7919) <= not((layer0_outputs(726)) or (layer0_outputs(7295)));
    layer1_outputs(7920) <= layer0_outputs(1218);
    layer1_outputs(7921) <= '0';
    layer1_outputs(7922) <= layer0_outputs(1743);
    layer1_outputs(7923) <= not(layer0_outputs(4120)) or (layer0_outputs(6796));
    layer1_outputs(7924) <= (layer0_outputs(9065)) xor (layer0_outputs(4112));
    layer1_outputs(7925) <= '0';
    layer1_outputs(7926) <= layer0_outputs(1641);
    layer1_outputs(7927) <= not(layer0_outputs(3729));
    layer1_outputs(7928) <= '0';
    layer1_outputs(7929) <= layer0_outputs(4188);
    layer1_outputs(7930) <= (layer0_outputs(2611)) xor (layer0_outputs(2274));
    layer1_outputs(7931) <= not(layer0_outputs(288)) or (layer0_outputs(579));
    layer1_outputs(7932) <= not((layer0_outputs(9121)) or (layer0_outputs(9272)));
    layer1_outputs(7933) <= not((layer0_outputs(6370)) and (layer0_outputs(4636)));
    layer1_outputs(7934) <= not(layer0_outputs(3552));
    layer1_outputs(7935) <= (layer0_outputs(6736)) and not (layer0_outputs(4857));
    layer1_outputs(7936) <= not(layer0_outputs(8784)) or (layer0_outputs(5012));
    layer1_outputs(7937) <= not(layer0_outputs(1943));
    layer1_outputs(7938) <= layer0_outputs(3404);
    layer1_outputs(7939) <= (layer0_outputs(6896)) and not (layer0_outputs(8927));
    layer1_outputs(7940) <= (layer0_outputs(6751)) and not (layer0_outputs(159));
    layer1_outputs(7941) <= layer0_outputs(8168);
    layer1_outputs(7942) <= (layer0_outputs(2667)) xor (layer0_outputs(6721));
    layer1_outputs(7943) <= not((layer0_outputs(1488)) and (layer0_outputs(4540)));
    layer1_outputs(7944) <= not(layer0_outputs(3737));
    layer1_outputs(7945) <= not(layer0_outputs(4978)) or (layer0_outputs(693));
    layer1_outputs(7946) <= not(layer0_outputs(6680)) or (layer0_outputs(4309));
    layer1_outputs(7947) <= not(layer0_outputs(9739));
    layer1_outputs(7948) <= layer0_outputs(2649);
    layer1_outputs(7949) <= '0';
    layer1_outputs(7950) <= not(layer0_outputs(1610));
    layer1_outputs(7951) <= (layer0_outputs(6281)) xor (layer0_outputs(81));
    layer1_outputs(7952) <= layer0_outputs(4754);
    layer1_outputs(7953) <= layer0_outputs(918);
    layer1_outputs(7954) <= layer0_outputs(6327);
    layer1_outputs(7955) <= not(layer0_outputs(1881));
    layer1_outputs(7956) <= (layer0_outputs(8684)) and (layer0_outputs(1811));
    layer1_outputs(7957) <= (layer0_outputs(78)) and not (layer0_outputs(7781));
    layer1_outputs(7958) <= not(layer0_outputs(887));
    layer1_outputs(7959) <= not(layer0_outputs(10155));
    layer1_outputs(7960) <= not(layer0_outputs(2189));
    layer1_outputs(7961) <= not(layer0_outputs(7594)) or (layer0_outputs(4034));
    layer1_outputs(7962) <= layer0_outputs(8087);
    layer1_outputs(7963) <= not((layer0_outputs(2303)) and (layer0_outputs(3992)));
    layer1_outputs(7964) <= not(layer0_outputs(8502));
    layer1_outputs(7965) <= not((layer0_outputs(6401)) and (layer0_outputs(7643)));
    layer1_outputs(7966) <= not(layer0_outputs(5495));
    layer1_outputs(7967) <= layer0_outputs(10050);
    layer1_outputs(7968) <= not((layer0_outputs(780)) xor (layer0_outputs(3951)));
    layer1_outputs(7969) <= not((layer0_outputs(5837)) xor (layer0_outputs(5097)));
    layer1_outputs(7970) <= (layer0_outputs(6134)) and (layer0_outputs(6042));
    layer1_outputs(7971) <= (layer0_outputs(4055)) and not (layer0_outputs(1040));
    layer1_outputs(7972) <= layer0_outputs(2504);
    layer1_outputs(7973) <= not(layer0_outputs(795));
    layer1_outputs(7974) <= (layer0_outputs(3736)) xor (layer0_outputs(5681));
    layer1_outputs(7975) <= not(layer0_outputs(9368));
    layer1_outputs(7976) <= (layer0_outputs(5780)) and not (layer0_outputs(3938));
    layer1_outputs(7977) <= (layer0_outputs(4037)) and (layer0_outputs(2671));
    layer1_outputs(7978) <= not(layer0_outputs(10226));
    layer1_outputs(7979) <= (layer0_outputs(7570)) and not (layer0_outputs(6146));
    layer1_outputs(7980) <= (layer0_outputs(3467)) and not (layer0_outputs(2452));
    layer1_outputs(7981) <= (layer0_outputs(10108)) and not (layer0_outputs(7701));
    layer1_outputs(7982) <= (layer0_outputs(694)) and (layer0_outputs(951));
    layer1_outputs(7983) <= layer0_outputs(9377);
    layer1_outputs(7984) <= (layer0_outputs(7900)) and not (layer0_outputs(2495));
    layer1_outputs(7985) <= layer0_outputs(6077);
    layer1_outputs(7986) <= (layer0_outputs(3056)) and not (layer0_outputs(709));
    layer1_outputs(7987) <= not((layer0_outputs(6324)) or (layer0_outputs(9274)));
    layer1_outputs(7988) <= layer0_outputs(3791);
    layer1_outputs(7989) <= not(layer0_outputs(4753));
    layer1_outputs(7990) <= not(layer0_outputs(2020));
    layer1_outputs(7991) <= layer0_outputs(8334);
    layer1_outputs(7992) <= not(layer0_outputs(8846)) or (layer0_outputs(5750));
    layer1_outputs(7993) <= not(layer0_outputs(8250));
    layer1_outputs(7994) <= not(layer0_outputs(9579));
    layer1_outputs(7995) <= (layer0_outputs(395)) and (layer0_outputs(10180));
    layer1_outputs(7996) <= not(layer0_outputs(2906));
    layer1_outputs(7997) <= not((layer0_outputs(5326)) or (layer0_outputs(1042)));
    layer1_outputs(7998) <= (layer0_outputs(8133)) and (layer0_outputs(4237));
    layer1_outputs(7999) <= not(layer0_outputs(3745));
    layer1_outputs(8000) <= (layer0_outputs(7513)) and not (layer0_outputs(10177));
    layer1_outputs(8001) <= layer0_outputs(2125);
    layer1_outputs(8002) <= not((layer0_outputs(4769)) or (layer0_outputs(5706)));
    layer1_outputs(8003) <= not(layer0_outputs(9096));
    layer1_outputs(8004) <= layer0_outputs(2143);
    layer1_outputs(8005) <= (layer0_outputs(2091)) and not (layer0_outputs(8491));
    layer1_outputs(8006) <= not((layer0_outputs(8139)) or (layer0_outputs(53)));
    layer1_outputs(8007) <= (layer0_outputs(7331)) and not (layer0_outputs(9503));
    layer1_outputs(8008) <= '0';
    layer1_outputs(8009) <= not(layer0_outputs(4570)) or (layer0_outputs(5074));
    layer1_outputs(8010) <= (layer0_outputs(7066)) and not (layer0_outputs(5143));
    layer1_outputs(8011) <= not((layer0_outputs(8801)) xor (layer0_outputs(86)));
    layer1_outputs(8012) <= (layer0_outputs(9256)) and not (layer0_outputs(5948));
    layer1_outputs(8013) <= not(layer0_outputs(8294)) or (layer0_outputs(6772));
    layer1_outputs(8014) <= (layer0_outputs(4801)) or (layer0_outputs(1847));
    layer1_outputs(8015) <= layer0_outputs(5390);
    layer1_outputs(8016) <= not(layer0_outputs(2452));
    layer1_outputs(8017) <= not(layer0_outputs(8886)) or (layer0_outputs(8098));
    layer1_outputs(8018) <= layer0_outputs(10226);
    layer1_outputs(8019) <= not(layer0_outputs(4634));
    layer1_outputs(8020) <= not(layer0_outputs(7141)) or (layer0_outputs(7930));
    layer1_outputs(8021) <= (layer0_outputs(8559)) or (layer0_outputs(3652));
    layer1_outputs(8022) <= '1';
    layer1_outputs(8023) <= not(layer0_outputs(2930));
    layer1_outputs(8024) <= (layer0_outputs(6058)) or (layer0_outputs(2630));
    layer1_outputs(8025) <= not(layer0_outputs(9825)) or (layer0_outputs(9094));
    layer1_outputs(8026) <= layer0_outputs(4335);
    layer1_outputs(8027) <= not(layer0_outputs(2170));
    layer1_outputs(8028) <= not(layer0_outputs(1489));
    layer1_outputs(8029) <= (layer0_outputs(8934)) and not (layer0_outputs(9419));
    layer1_outputs(8030) <= not((layer0_outputs(7786)) xor (layer0_outputs(1707)));
    layer1_outputs(8031) <= not(layer0_outputs(4911)) or (layer0_outputs(5631));
    layer1_outputs(8032) <= not((layer0_outputs(451)) and (layer0_outputs(6433)));
    layer1_outputs(8033) <= not((layer0_outputs(5387)) or (layer0_outputs(5312)));
    layer1_outputs(8034) <= not((layer0_outputs(7365)) xor (layer0_outputs(3924)));
    layer1_outputs(8035) <= (layer0_outputs(5222)) and not (layer0_outputs(7546));
    layer1_outputs(8036) <= '1';
    layer1_outputs(8037) <= layer0_outputs(8326);
    layer1_outputs(8038) <= (layer0_outputs(9544)) and not (layer0_outputs(6153));
    layer1_outputs(8039) <= not((layer0_outputs(6615)) xor (layer0_outputs(2685)));
    layer1_outputs(8040) <= not(layer0_outputs(3818));
    layer1_outputs(8041) <= (layer0_outputs(2698)) or (layer0_outputs(1629));
    layer1_outputs(8042) <= layer0_outputs(2801);
    layer1_outputs(8043) <= (layer0_outputs(9751)) or (layer0_outputs(6785));
    layer1_outputs(8044) <= (layer0_outputs(6829)) and not (layer0_outputs(1182));
    layer1_outputs(8045) <= not(layer0_outputs(6734));
    layer1_outputs(8046) <= (layer0_outputs(10148)) and not (layer0_outputs(7136));
    layer1_outputs(8047) <= not((layer0_outputs(4759)) or (layer0_outputs(3240)));
    layer1_outputs(8048) <= not(layer0_outputs(5200));
    layer1_outputs(8049) <= (layer0_outputs(1668)) or (layer0_outputs(5958));
    layer1_outputs(8050) <= '0';
    layer1_outputs(8051) <= layer0_outputs(7882);
    layer1_outputs(8052) <= not((layer0_outputs(5676)) or (layer0_outputs(1344)));
    layer1_outputs(8053) <= not(layer0_outputs(10021));
    layer1_outputs(8054) <= layer0_outputs(3378);
    layer1_outputs(8055) <= not((layer0_outputs(1193)) xor (layer0_outputs(7714)));
    layer1_outputs(8056) <= not(layer0_outputs(3046));
    layer1_outputs(8057) <= (layer0_outputs(3977)) and not (layer0_outputs(1928));
    layer1_outputs(8058) <= layer0_outputs(8691);
    layer1_outputs(8059) <= not(layer0_outputs(8286));
    layer1_outputs(8060) <= '1';
    layer1_outputs(8061) <= (layer0_outputs(5242)) and not (layer0_outputs(1346));
    layer1_outputs(8062) <= (layer0_outputs(5366)) and not (layer0_outputs(2078));
    layer1_outputs(8063) <= '1';
    layer1_outputs(8064) <= layer0_outputs(8590);
    layer1_outputs(8065) <= (layer0_outputs(9530)) and (layer0_outputs(6813));
    layer1_outputs(8066) <= (layer0_outputs(8503)) and (layer0_outputs(3214));
    layer1_outputs(8067) <= (layer0_outputs(6662)) and not (layer0_outputs(1004));
    layer1_outputs(8068) <= not(layer0_outputs(635)) or (layer0_outputs(810));
    layer1_outputs(8069) <= not(layer0_outputs(9348));
    layer1_outputs(8070) <= (layer0_outputs(2405)) or (layer0_outputs(1270));
    layer1_outputs(8071) <= not(layer0_outputs(304));
    layer1_outputs(8072) <= not(layer0_outputs(2919)) or (layer0_outputs(2900));
    layer1_outputs(8073) <= not((layer0_outputs(6893)) xor (layer0_outputs(8846)));
    layer1_outputs(8074) <= (layer0_outputs(1744)) and (layer0_outputs(7747));
    layer1_outputs(8075) <= layer0_outputs(3101);
    layer1_outputs(8076) <= not((layer0_outputs(2188)) or (layer0_outputs(9758)));
    layer1_outputs(8077) <= not(layer0_outputs(4004)) or (layer0_outputs(112));
    layer1_outputs(8078) <= (layer0_outputs(3886)) xor (layer0_outputs(4696));
    layer1_outputs(8079) <= layer0_outputs(3869);
    layer1_outputs(8080) <= not(layer0_outputs(3289));
    layer1_outputs(8081) <= not(layer0_outputs(2734)) or (layer0_outputs(10231));
    layer1_outputs(8082) <= (layer0_outputs(1171)) and not (layer0_outputs(9273));
    layer1_outputs(8083) <= layer0_outputs(7683);
    layer1_outputs(8084) <= not((layer0_outputs(7802)) or (layer0_outputs(8919)));
    layer1_outputs(8085) <= '0';
    layer1_outputs(8086) <= not((layer0_outputs(9016)) and (layer0_outputs(5159)));
    layer1_outputs(8087) <= (layer0_outputs(3504)) and not (layer0_outputs(3222));
    layer1_outputs(8088) <= not(layer0_outputs(4235));
    layer1_outputs(8089) <= not(layer0_outputs(10043));
    layer1_outputs(8090) <= not(layer0_outputs(2476));
    layer1_outputs(8091) <= not((layer0_outputs(1648)) and (layer0_outputs(7980)));
    layer1_outputs(8092) <= layer0_outputs(1661);
    layer1_outputs(8093) <= layer0_outputs(7123);
    layer1_outputs(8094) <= not(layer0_outputs(9079));
    layer1_outputs(8095) <= (layer0_outputs(7692)) xor (layer0_outputs(3535));
    layer1_outputs(8096) <= not(layer0_outputs(7061));
    layer1_outputs(8097) <= not(layer0_outputs(850));
    layer1_outputs(8098) <= layer0_outputs(6474);
    layer1_outputs(8099) <= not(layer0_outputs(3945));
    layer1_outputs(8100) <= not(layer0_outputs(7438));
    layer1_outputs(8101) <= not(layer0_outputs(4694)) or (layer0_outputs(8682));
    layer1_outputs(8102) <= layer0_outputs(5606);
    layer1_outputs(8103) <= not(layer0_outputs(4729)) or (layer0_outputs(6070));
    layer1_outputs(8104) <= (layer0_outputs(9681)) and (layer0_outputs(4311));
    layer1_outputs(8105) <= not((layer0_outputs(9312)) or (layer0_outputs(9046)));
    layer1_outputs(8106) <= not(layer0_outputs(5322));
    layer1_outputs(8107) <= not(layer0_outputs(19)) or (layer0_outputs(6873));
    layer1_outputs(8108) <= (layer0_outputs(7374)) and not (layer0_outputs(8160));
    layer1_outputs(8109) <= not(layer0_outputs(2560));
    layer1_outputs(8110) <= not(layer0_outputs(9318));
    layer1_outputs(8111) <= not(layer0_outputs(2607));
    layer1_outputs(8112) <= layer0_outputs(7281);
    layer1_outputs(8113) <= not((layer0_outputs(6556)) and (layer0_outputs(2908)));
    layer1_outputs(8114) <= not(layer0_outputs(2020));
    layer1_outputs(8115) <= not(layer0_outputs(3672)) or (layer0_outputs(9710));
    layer1_outputs(8116) <= (layer0_outputs(8791)) or (layer0_outputs(9239));
    layer1_outputs(8117) <= not(layer0_outputs(7234));
    layer1_outputs(8118) <= layer0_outputs(3802);
    layer1_outputs(8119) <= not(layer0_outputs(7816));
    layer1_outputs(8120) <= (layer0_outputs(901)) and not (layer0_outputs(5507));
    layer1_outputs(8121) <= (layer0_outputs(5461)) xor (layer0_outputs(5205));
    layer1_outputs(8122) <= (layer0_outputs(6881)) or (layer0_outputs(7503));
    layer1_outputs(8123) <= layer0_outputs(8114);
    layer1_outputs(8124) <= not((layer0_outputs(937)) or (layer0_outputs(128)));
    layer1_outputs(8125) <= '0';
    layer1_outputs(8126) <= '0';
    layer1_outputs(8127) <= not(layer0_outputs(3824)) or (layer0_outputs(2428));
    layer1_outputs(8128) <= not((layer0_outputs(1327)) xor (layer0_outputs(846)));
    layer1_outputs(8129) <= not(layer0_outputs(3747)) or (layer0_outputs(5519));
    layer1_outputs(8130) <= not(layer0_outputs(6657));
    layer1_outputs(8131) <= not(layer0_outputs(7222));
    layer1_outputs(8132) <= (layer0_outputs(1354)) and (layer0_outputs(2551));
    layer1_outputs(8133) <= not((layer0_outputs(8661)) or (layer0_outputs(5740)));
    layer1_outputs(8134) <= layer0_outputs(5414);
    layer1_outputs(8135) <= (layer0_outputs(785)) and not (layer0_outputs(751));
    layer1_outputs(8136) <= not(layer0_outputs(1822));
    layer1_outputs(8137) <= layer0_outputs(5361);
    layer1_outputs(8138) <= not(layer0_outputs(2154)) or (layer0_outputs(4150));
    layer1_outputs(8139) <= (layer0_outputs(9522)) and not (layer0_outputs(3432));
    layer1_outputs(8140) <= not((layer0_outputs(5922)) or (layer0_outputs(4945)));
    layer1_outputs(8141) <= not((layer0_outputs(3989)) xor (layer0_outputs(5121)));
    layer1_outputs(8142) <= '0';
    layer1_outputs(8143) <= (layer0_outputs(6038)) or (layer0_outputs(3605));
    layer1_outputs(8144) <= not(layer0_outputs(1885)) or (layer0_outputs(9456));
    layer1_outputs(8145) <= not(layer0_outputs(7323));
    layer1_outputs(8146) <= not(layer0_outputs(4024)) or (layer0_outputs(1257));
    layer1_outputs(8147) <= not(layer0_outputs(4823));
    layer1_outputs(8148) <= (layer0_outputs(7148)) xor (layer0_outputs(1205));
    layer1_outputs(8149) <= layer0_outputs(9039);
    layer1_outputs(8150) <= layer0_outputs(4640);
    layer1_outputs(8151) <= not((layer0_outputs(1630)) or (layer0_outputs(7886)));
    layer1_outputs(8152) <= layer0_outputs(2549);
    layer1_outputs(8153) <= layer0_outputs(1337);
    layer1_outputs(8154) <= not(layer0_outputs(8041)) or (layer0_outputs(10132));
    layer1_outputs(8155) <= not(layer0_outputs(2223));
    layer1_outputs(8156) <= (layer0_outputs(8396)) and (layer0_outputs(3389));
    layer1_outputs(8157) <= (layer0_outputs(7349)) xor (layer0_outputs(8458));
    layer1_outputs(8158) <= '1';
    layer1_outputs(8159) <= (layer0_outputs(6907)) xor (layer0_outputs(6384));
    layer1_outputs(8160) <= (layer0_outputs(1559)) xor (layer0_outputs(5675));
    layer1_outputs(8161) <= layer0_outputs(2058);
    layer1_outputs(8162) <= not((layer0_outputs(4416)) xor (layer0_outputs(9505)));
    layer1_outputs(8163) <= layer0_outputs(6101);
    layer1_outputs(8164) <= (layer0_outputs(3217)) and not (layer0_outputs(8608));
    layer1_outputs(8165) <= (layer0_outputs(2236)) or (layer0_outputs(5117));
    layer1_outputs(8166) <= (layer0_outputs(6571)) and not (layer0_outputs(1986));
    layer1_outputs(8167) <= not(layer0_outputs(477));
    layer1_outputs(8168) <= (layer0_outputs(7904)) or (layer0_outputs(8881));
    layer1_outputs(8169) <= not(layer0_outputs(6404));
    layer1_outputs(8170) <= not((layer0_outputs(9847)) and (layer0_outputs(7042)));
    layer1_outputs(8171) <= layer0_outputs(9754);
    layer1_outputs(8172) <= not(layer0_outputs(4437));
    layer1_outputs(8173) <= layer0_outputs(2286);
    layer1_outputs(8174) <= not(layer0_outputs(1045)) or (layer0_outputs(8751));
    layer1_outputs(8175) <= not(layer0_outputs(937));
    layer1_outputs(8176) <= not(layer0_outputs(1791)) or (layer0_outputs(7557));
    layer1_outputs(8177) <= '0';
    layer1_outputs(8178) <= not(layer0_outputs(4529));
    layer1_outputs(8179) <= (layer0_outputs(853)) or (layer0_outputs(10229));
    layer1_outputs(8180) <= not((layer0_outputs(2528)) or (layer0_outputs(9880)));
    layer1_outputs(8181) <= '0';
    layer1_outputs(8182) <= not(layer0_outputs(4593));
    layer1_outputs(8183) <= not(layer0_outputs(9042)) or (layer0_outputs(1329));
    layer1_outputs(8184) <= not((layer0_outputs(3814)) or (layer0_outputs(4476)));
    layer1_outputs(8185) <= '0';
    layer1_outputs(8186) <= not(layer0_outputs(605));
    layer1_outputs(8187) <= not((layer0_outputs(9925)) or (layer0_outputs(1955)));
    layer1_outputs(8188) <= not(layer0_outputs(1744));
    layer1_outputs(8189) <= (layer0_outputs(2086)) xor (layer0_outputs(1944));
    layer1_outputs(8190) <= layer0_outputs(5141);
    layer1_outputs(8191) <= not(layer0_outputs(7631));
    layer1_outputs(8192) <= layer0_outputs(7065);
    layer1_outputs(8193) <= not(layer0_outputs(83));
    layer1_outputs(8194) <= (layer0_outputs(5861)) and not (layer0_outputs(4430));
    layer1_outputs(8195) <= not(layer0_outputs(757)) or (layer0_outputs(209));
    layer1_outputs(8196) <= (layer0_outputs(6477)) or (layer0_outputs(5415));
    layer1_outputs(8197) <= not(layer0_outputs(3874)) or (layer0_outputs(9483));
    layer1_outputs(8198) <= layer0_outputs(3484);
    layer1_outputs(8199) <= '0';
    layer1_outputs(8200) <= (layer0_outputs(1376)) or (layer0_outputs(6279));
    layer1_outputs(8201) <= not((layer0_outputs(7436)) and (layer0_outputs(7206)));
    layer1_outputs(8202) <= not(layer0_outputs(2828)) or (layer0_outputs(10066));
    layer1_outputs(8203) <= (layer0_outputs(8708)) and not (layer0_outputs(9182));
    layer1_outputs(8204) <= not((layer0_outputs(8125)) or (layer0_outputs(2935)));
    layer1_outputs(8205) <= not((layer0_outputs(1851)) or (layer0_outputs(702)));
    layer1_outputs(8206) <= (layer0_outputs(1349)) and not (layer0_outputs(9434));
    layer1_outputs(8207) <= layer0_outputs(6080);
    layer1_outputs(8208) <= not(layer0_outputs(1355)) or (layer0_outputs(962));
    layer1_outputs(8209) <= layer0_outputs(7082);
    layer1_outputs(8210) <= not(layer0_outputs(6765));
    layer1_outputs(8211) <= not(layer0_outputs(5335)) or (layer0_outputs(7037));
    layer1_outputs(8212) <= layer0_outputs(6918);
    layer1_outputs(8213) <= not((layer0_outputs(8765)) and (layer0_outputs(1404)));
    layer1_outputs(8214) <= not((layer0_outputs(556)) xor (layer0_outputs(6858)));
    layer1_outputs(8215) <= (layer0_outputs(6206)) or (layer0_outputs(7298));
    layer1_outputs(8216) <= layer0_outputs(3916);
    layer1_outputs(8217) <= not(layer0_outputs(7626));
    layer1_outputs(8218) <= (layer0_outputs(1732)) xor (layer0_outputs(2334));
    layer1_outputs(8219) <= not((layer0_outputs(827)) or (layer0_outputs(3947)));
    layer1_outputs(8220) <= not(layer0_outputs(7220));
    layer1_outputs(8221) <= not(layer0_outputs(6820));
    layer1_outputs(8222) <= not(layer0_outputs(151)) or (layer0_outputs(2920));
    layer1_outputs(8223) <= not((layer0_outputs(7207)) and (layer0_outputs(981)));
    layer1_outputs(8224) <= not(layer0_outputs(5448)) or (layer0_outputs(1834));
    layer1_outputs(8225) <= layer0_outputs(5982);
    layer1_outputs(8226) <= (layer0_outputs(1056)) and not (layer0_outputs(891));
    layer1_outputs(8227) <= not(layer0_outputs(5335));
    layer1_outputs(8228) <= (layer0_outputs(1313)) and (layer0_outputs(3933));
    layer1_outputs(8229) <= (layer0_outputs(1463)) or (layer0_outputs(5745));
    layer1_outputs(8230) <= (layer0_outputs(6812)) and not (layer0_outputs(10230));
    layer1_outputs(8231) <= (layer0_outputs(3718)) xor (layer0_outputs(9299));
    layer1_outputs(8232) <= not(layer0_outputs(6976)) or (layer0_outputs(3155));
    layer1_outputs(8233) <= not(layer0_outputs(5205));
    layer1_outputs(8234) <= not(layer0_outputs(4113));
    layer1_outputs(8235) <= (layer0_outputs(9684)) and not (layer0_outputs(2467));
    layer1_outputs(8236) <= (layer0_outputs(1293)) and not (layer0_outputs(3837));
    layer1_outputs(8237) <= not(layer0_outputs(7535));
    layer1_outputs(8238) <= not(layer0_outputs(2790));
    layer1_outputs(8239) <= not(layer0_outputs(4018));
    layer1_outputs(8240) <= layer0_outputs(2204);
    layer1_outputs(8241) <= (layer0_outputs(9658)) and not (layer0_outputs(6154));
    layer1_outputs(8242) <= layer0_outputs(6693);
    layer1_outputs(8243) <= layer0_outputs(955);
    layer1_outputs(8244) <= not(layer0_outputs(9220));
    layer1_outputs(8245) <= '0';
    layer1_outputs(8246) <= layer0_outputs(8642);
    layer1_outputs(8247) <= (layer0_outputs(1334)) and (layer0_outputs(3253));
    layer1_outputs(8248) <= (layer0_outputs(2416)) and (layer0_outputs(4325));
    layer1_outputs(8249) <= not(layer0_outputs(5574));
    layer1_outputs(8250) <= (layer0_outputs(2454)) or (layer0_outputs(8442));
    layer1_outputs(8251) <= not((layer0_outputs(9484)) or (layer0_outputs(8110)));
    layer1_outputs(8252) <= '0';
    layer1_outputs(8253) <= not(layer0_outputs(5526)) or (layer0_outputs(1268));
    layer1_outputs(8254) <= (layer0_outputs(1494)) and not (layer0_outputs(201));
    layer1_outputs(8255) <= (layer0_outputs(8643)) or (layer0_outputs(8976));
    layer1_outputs(8256) <= not(layer0_outputs(622));
    layer1_outputs(8257) <= '0';
    layer1_outputs(8258) <= not(layer0_outputs(3489));
    layer1_outputs(8259) <= (layer0_outputs(7055)) or (layer0_outputs(8955));
    layer1_outputs(8260) <= not(layer0_outputs(2779));
    layer1_outputs(8261) <= not(layer0_outputs(8645)) or (layer0_outputs(1681));
    layer1_outputs(8262) <= not(layer0_outputs(2657));
    layer1_outputs(8263) <= (layer0_outputs(6287)) and not (layer0_outputs(5438));
    layer1_outputs(8264) <= not(layer0_outputs(6946)) or (layer0_outputs(7686));
    layer1_outputs(8265) <= (layer0_outputs(5434)) and (layer0_outputs(8483));
    layer1_outputs(8266) <= (layer0_outputs(5449)) and not (layer0_outputs(7837));
    layer1_outputs(8267) <= '0';
    layer1_outputs(8268) <= not(layer0_outputs(7174));
    layer1_outputs(8269) <= not(layer0_outputs(7077));
    layer1_outputs(8270) <= not((layer0_outputs(7499)) and (layer0_outputs(129)));
    layer1_outputs(8271) <= layer0_outputs(9814);
    layer1_outputs(8272) <= not((layer0_outputs(2164)) xor (layer0_outputs(3003)));
    layer1_outputs(8273) <= not(layer0_outputs(7907));
    layer1_outputs(8274) <= not((layer0_outputs(8911)) and (layer0_outputs(7434)));
    layer1_outputs(8275) <= layer0_outputs(4820);
    layer1_outputs(8276) <= not(layer0_outputs(10090)) or (layer0_outputs(9683));
    layer1_outputs(8277) <= (layer0_outputs(8646)) and (layer0_outputs(9642));
    layer1_outputs(8278) <= (layer0_outputs(743)) and not (layer0_outputs(3485));
    layer1_outputs(8279) <= (layer0_outputs(1867)) or (layer0_outputs(7906));
    layer1_outputs(8280) <= (layer0_outputs(442)) or (layer0_outputs(3022));
    layer1_outputs(8281) <= not(layer0_outputs(4665)) or (layer0_outputs(2658));
    layer1_outputs(8282) <= not((layer0_outputs(1196)) and (layer0_outputs(4295)));
    layer1_outputs(8283) <= not(layer0_outputs(5128));
    layer1_outputs(8284) <= not(layer0_outputs(5091)) or (layer0_outputs(5755));
    layer1_outputs(8285) <= not((layer0_outputs(1779)) and (layer0_outputs(950)));
    layer1_outputs(8286) <= (layer0_outputs(3190)) and (layer0_outputs(5306));
    layer1_outputs(8287) <= '0';
    layer1_outputs(8288) <= not((layer0_outputs(1601)) or (layer0_outputs(9020)));
    layer1_outputs(8289) <= not((layer0_outputs(2276)) and (layer0_outputs(1800)));
    layer1_outputs(8290) <= not(layer0_outputs(3725)) or (layer0_outputs(3879));
    layer1_outputs(8291) <= not((layer0_outputs(3248)) xor (layer0_outputs(9296)));
    layer1_outputs(8292) <= not((layer0_outputs(9704)) xor (layer0_outputs(6853)));
    layer1_outputs(8293) <= layer0_outputs(7699);
    layer1_outputs(8294) <= not((layer0_outputs(8531)) and (layer0_outputs(7476)));
    layer1_outputs(8295) <= (layer0_outputs(2168)) or (layer0_outputs(315));
    layer1_outputs(8296) <= not(layer0_outputs(44));
    layer1_outputs(8297) <= layer0_outputs(783);
    layer1_outputs(8298) <= (layer0_outputs(10136)) and (layer0_outputs(2441));
    layer1_outputs(8299) <= not(layer0_outputs(4466));
    layer1_outputs(8300) <= (layer0_outputs(10137)) and (layer0_outputs(8079));
    layer1_outputs(8301) <= (layer0_outputs(8021)) and not (layer0_outputs(6072));
    layer1_outputs(8302) <= '1';
    layer1_outputs(8303) <= not(layer0_outputs(444)) or (layer0_outputs(1375));
    layer1_outputs(8304) <= (layer0_outputs(5360)) xor (layer0_outputs(4681));
    layer1_outputs(8305) <= layer0_outputs(6706);
    layer1_outputs(8306) <= not(layer0_outputs(1360));
    layer1_outputs(8307) <= (layer0_outputs(8810)) and (layer0_outputs(8077));
    layer1_outputs(8308) <= (layer0_outputs(7958)) and not (layer0_outputs(999));
    layer1_outputs(8309) <= (layer0_outputs(1315)) xor (layer0_outputs(3870));
    layer1_outputs(8310) <= (layer0_outputs(4734)) xor (layer0_outputs(7276));
    layer1_outputs(8311) <= layer0_outputs(6364);
    layer1_outputs(8312) <= not((layer0_outputs(8211)) and (layer0_outputs(1155)));
    layer1_outputs(8313) <= not(layer0_outputs(6583)) or (layer0_outputs(1448));
    layer1_outputs(8314) <= not(layer0_outputs(2417));
    layer1_outputs(8315) <= (layer0_outputs(3426)) and not (layer0_outputs(10105));
    layer1_outputs(8316) <= (layer0_outputs(8470)) and not (layer0_outputs(5456));
    layer1_outputs(8317) <= not(layer0_outputs(6377)) or (layer0_outputs(2257));
    layer1_outputs(8318) <= (layer0_outputs(9823)) and (layer0_outputs(3308));
    layer1_outputs(8319) <= (layer0_outputs(5512)) or (layer0_outputs(187));
    layer1_outputs(8320) <= not(layer0_outputs(2614));
    layer1_outputs(8321) <= (layer0_outputs(6649)) xor (layer0_outputs(5846));
    layer1_outputs(8322) <= not((layer0_outputs(3437)) and (layer0_outputs(4245)));
    layer1_outputs(8323) <= not((layer0_outputs(6149)) and (layer0_outputs(5920)));
    layer1_outputs(8324) <= not(layer0_outputs(10068));
    layer1_outputs(8325) <= layer0_outputs(9184);
    layer1_outputs(8326) <= '0';
    layer1_outputs(8327) <= (layer0_outputs(2034)) and not (layer0_outputs(8396));
    layer1_outputs(8328) <= (layer0_outputs(3817)) and not (layer0_outputs(1887));
    layer1_outputs(8329) <= layer0_outputs(6235);
    layer1_outputs(8330) <= layer0_outputs(5887);
    layer1_outputs(8331) <= layer0_outputs(7737);
    layer1_outputs(8332) <= '1';
    layer1_outputs(8333) <= not((layer0_outputs(3477)) xor (layer0_outputs(7573)));
    layer1_outputs(8334) <= (layer0_outputs(8006)) or (layer0_outputs(7074));
    layer1_outputs(8335) <= (layer0_outputs(3607)) or (layer0_outputs(3475));
    layer1_outputs(8336) <= '1';
    layer1_outputs(8337) <= not(layer0_outputs(1054));
    layer1_outputs(8338) <= not(layer0_outputs(8720)) or (layer0_outputs(3843));
    layer1_outputs(8339) <= layer0_outputs(8552);
    layer1_outputs(8340) <= not(layer0_outputs(6954)) or (layer0_outputs(9296));
    layer1_outputs(8341) <= not(layer0_outputs(4882));
    layer1_outputs(8342) <= layer0_outputs(7655);
    layer1_outputs(8343) <= (layer0_outputs(6750)) and (layer0_outputs(1451));
    layer1_outputs(8344) <= not(layer0_outputs(124));
    layer1_outputs(8345) <= not(layer0_outputs(1692)) or (layer0_outputs(9607));
    layer1_outputs(8346) <= (layer0_outputs(10032)) or (layer0_outputs(1285));
    layer1_outputs(8347) <= not(layer0_outputs(7220));
    layer1_outputs(8348) <= not(layer0_outputs(7558));
    layer1_outputs(8349) <= not(layer0_outputs(1456));
    layer1_outputs(8350) <= not((layer0_outputs(1984)) xor (layer0_outputs(6238)));
    layer1_outputs(8351) <= (layer0_outputs(1609)) and not (layer0_outputs(2835));
    layer1_outputs(8352) <= layer0_outputs(3834);
    layer1_outputs(8353) <= not((layer0_outputs(8961)) xor (layer0_outputs(1257)));
    layer1_outputs(8354) <= layer0_outputs(9755);
    layer1_outputs(8355) <= not(layer0_outputs(1277)) or (layer0_outputs(6409));
    layer1_outputs(8356) <= not((layer0_outputs(9898)) or (layer0_outputs(5698)));
    layer1_outputs(8357) <= layer0_outputs(2871);
    layer1_outputs(8358) <= not(layer0_outputs(2923));
    layer1_outputs(8359) <= layer0_outputs(837);
    layer1_outputs(8360) <= layer0_outputs(1597);
    layer1_outputs(8361) <= not((layer0_outputs(2109)) or (layer0_outputs(2357)));
    layer1_outputs(8362) <= layer0_outputs(7659);
    layer1_outputs(8363) <= layer0_outputs(7443);
    layer1_outputs(8364) <= (layer0_outputs(3942)) and (layer0_outputs(9619));
    layer1_outputs(8365) <= not(layer0_outputs(10065)) or (layer0_outputs(875));
    layer1_outputs(8366) <= not(layer0_outputs(3863));
    layer1_outputs(8367) <= (layer0_outputs(4975)) and not (layer0_outputs(4762));
    layer1_outputs(8368) <= not((layer0_outputs(3843)) or (layer0_outputs(6120)));
    layer1_outputs(8369) <= (layer0_outputs(4569)) xor (layer0_outputs(5586));
    layer1_outputs(8370) <= not((layer0_outputs(4088)) or (layer0_outputs(707)));
    layer1_outputs(8371) <= not(layer0_outputs(9612));
    layer1_outputs(8372) <= not(layer0_outputs(7976)) or (layer0_outputs(2333));
    layer1_outputs(8373) <= (layer0_outputs(6432)) and (layer0_outputs(7500));
    layer1_outputs(8374) <= not((layer0_outputs(5063)) or (layer0_outputs(4666)));
    layer1_outputs(8375) <= not(layer0_outputs(6141)) or (layer0_outputs(6024));
    layer1_outputs(8376) <= not((layer0_outputs(7497)) or (layer0_outputs(9797)));
    layer1_outputs(8377) <= not(layer0_outputs(2665)) or (layer0_outputs(9911));
    layer1_outputs(8378) <= '1';
    layer1_outputs(8379) <= not(layer0_outputs(8855)) or (layer0_outputs(3663));
    layer1_outputs(8380) <= layer0_outputs(6823);
    layer1_outputs(8381) <= not(layer0_outputs(3724)) or (layer0_outputs(5453));
    layer1_outputs(8382) <= not(layer0_outputs(8318));
    layer1_outputs(8383) <= not((layer0_outputs(6190)) or (layer0_outputs(7949)));
    layer1_outputs(8384) <= layer0_outputs(5644);
    layer1_outputs(8385) <= (layer0_outputs(8252)) and (layer0_outputs(10237));
    layer1_outputs(8386) <= not((layer0_outputs(6268)) xor (layer0_outputs(1777)));
    layer1_outputs(8387) <= layer0_outputs(1232);
    layer1_outputs(8388) <= '0';
    layer1_outputs(8389) <= (layer0_outputs(8601)) and (layer0_outputs(173));
    layer1_outputs(8390) <= (layer0_outputs(2227)) xor (layer0_outputs(1255));
    layer1_outputs(8391) <= (layer0_outputs(5158)) or (layer0_outputs(8742));
    layer1_outputs(8392) <= '0';
    layer1_outputs(8393) <= not(layer0_outputs(3696)) or (layer0_outputs(8359));
    layer1_outputs(8394) <= (layer0_outputs(7492)) or (layer0_outputs(4541));
    layer1_outputs(8395) <= (layer0_outputs(9610)) and (layer0_outputs(9877));
    layer1_outputs(8396) <= not((layer0_outputs(8174)) or (layer0_outputs(597)));
    layer1_outputs(8397) <= layer0_outputs(607);
    layer1_outputs(8398) <= layer0_outputs(8758);
    layer1_outputs(8399) <= not(layer0_outputs(3167)) or (layer0_outputs(9272));
    layer1_outputs(8400) <= layer0_outputs(7218);
    layer1_outputs(8401) <= not(layer0_outputs(3343));
    layer1_outputs(8402) <= not((layer0_outputs(5841)) and (layer0_outputs(4927)));
    layer1_outputs(8403) <= (layer0_outputs(6275)) and (layer0_outputs(1937));
    layer1_outputs(8404) <= layer0_outputs(9093);
    layer1_outputs(8405) <= not(layer0_outputs(9459));
    layer1_outputs(8406) <= not(layer0_outputs(8795));
    layer1_outputs(8407) <= not((layer0_outputs(3354)) xor (layer0_outputs(8500)));
    layer1_outputs(8408) <= not(layer0_outputs(1677)) or (layer0_outputs(3442));
    layer1_outputs(8409) <= layer0_outputs(8874);
    layer1_outputs(8410) <= not(layer0_outputs(3569));
    layer1_outputs(8411) <= not((layer0_outputs(2076)) or (layer0_outputs(9692)));
    layer1_outputs(8412) <= (layer0_outputs(6601)) and (layer0_outputs(4164));
    layer1_outputs(8413) <= (layer0_outputs(2207)) and (layer0_outputs(5710));
    layer1_outputs(8414) <= not(layer0_outputs(7685));
    layer1_outputs(8415) <= not(layer0_outputs(8465)) or (layer0_outputs(7348));
    layer1_outputs(8416) <= not((layer0_outputs(7463)) or (layer0_outputs(893)));
    layer1_outputs(8417) <= layer0_outputs(1075);
    layer1_outputs(8418) <= (layer0_outputs(5407)) and not (layer0_outputs(7646));
    layer1_outputs(8419) <= layer0_outputs(4506);
    layer1_outputs(8420) <= not((layer0_outputs(4378)) xor (layer0_outputs(5538)));
    layer1_outputs(8421) <= (layer0_outputs(243)) xor (layer0_outputs(8425));
    layer1_outputs(8422) <= not((layer0_outputs(8815)) or (layer0_outputs(6890)));
    layer1_outputs(8423) <= (layer0_outputs(2273)) and not (layer0_outputs(9409));
    layer1_outputs(8424) <= layer0_outputs(1847);
    layer1_outputs(8425) <= not((layer0_outputs(5754)) xor (layer0_outputs(7452)));
    layer1_outputs(8426) <= layer0_outputs(1103);
    layer1_outputs(8427) <= layer0_outputs(8932);
    layer1_outputs(8428) <= (layer0_outputs(8131)) and not (layer0_outputs(146));
    layer1_outputs(8429) <= not((layer0_outputs(4518)) or (layer0_outputs(10049)));
    layer1_outputs(8430) <= layer0_outputs(6311);
    layer1_outputs(8431) <= (layer0_outputs(3973)) and not (layer0_outputs(8480));
    layer1_outputs(8432) <= layer0_outputs(6155);
    layer1_outputs(8433) <= (layer0_outputs(2561)) and (layer0_outputs(5470));
    layer1_outputs(8434) <= layer0_outputs(8920);
    layer1_outputs(8435) <= not((layer0_outputs(5679)) xor (layer0_outputs(780)));
    layer1_outputs(8436) <= not(layer0_outputs(7237));
    layer1_outputs(8437) <= (layer0_outputs(1606)) and not (layer0_outputs(8264));
    layer1_outputs(8438) <= not((layer0_outputs(791)) and (layer0_outputs(125)));
    layer1_outputs(8439) <= not((layer0_outputs(6239)) or (layer0_outputs(3731)));
    layer1_outputs(8440) <= not((layer0_outputs(5796)) xor (layer0_outputs(312)));
    layer1_outputs(8441) <= layer0_outputs(2988);
    layer1_outputs(8442) <= not(layer0_outputs(2589)) or (layer0_outputs(7426));
    layer1_outputs(8443) <= (layer0_outputs(2827)) and not (layer0_outputs(6566));
    layer1_outputs(8444) <= not(layer0_outputs(6722));
    layer1_outputs(8445) <= not((layer0_outputs(1565)) and (layer0_outputs(7700)));
    layer1_outputs(8446) <= (layer0_outputs(8304)) and not (layer0_outputs(1979));
    layer1_outputs(8447) <= not((layer0_outputs(5408)) or (layer0_outputs(7784)));
    layer1_outputs(8448) <= (layer0_outputs(4869)) or (layer0_outputs(3804));
    layer1_outputs(8449) <= not((layer0_outputs(7223)) or (layer0_outputs(7778)));
    layer1_outputs(8450) <= not(layer0_outputs(6359));
    layer1_outputs(8451) <= layer0_outputs(5935);
    layer1_outputs(8452) <= layer0_outputs(1879);
    layer1_outputs(8453) <= not((layer0_outputs(7556)) or (layer0_outputs(1691)));
    layer1_outputs(8454) <= not(layer0_outputs(1765));
    layer1_outputs(8455) <= not(layer0_outputs(5026));
    layer1_outputs(8456) <= not((layer0_outputs(2290)) xor (layer0_outputs(3930)));
    layer1_outputs(8457) <= layer0_outputs(3773);
    layer1_outputs(8458) <= not(layer0_outputs(421));
    layer1_outputs(8459) <= not((layer0_outputs(736)) xor (layer0_outputs(729)));
    layer1_outputs(8460) <= (layer0_outputs(2236)) and not (layer0_outputs(4501));
    layer1_outputs(8461) <= (layer0_outputs(4405)) and (layer0_outputs(1170));
    layer1_outputs(8462) <= layer0_outputs(6517);
    layer1_outputs(8463) <= not(layer0_outputs(3509));
    layer1_outputs(8464) <= layer0_outputs(4697);
    layer1_outputs(8465) <= (layer0_outputs(2597)) and not (layer0_outputs(387));
    layer1_outputs(8466) <= (layer0_outputs(8613)) xor (layer0_outputs(7013));
    layer1_outputs(8467) <= (layer0_outputs(2630)) and not (layer0_outputs(1511));
    layer1_outputs(8468) <= (layer0_outputs(1060)) and not (layer0_outputs(8253));
    layer1_outputs(8469) <= layer0_outputs(7316);
    layer1_outputs(8470) <= not(layer0_outputs(864));
    layer1_outputs(8471) <= not(layer0_outputs(136));
    layer1_outputs(8472) <= '1';
    layer1_outputs(8473) <= not(layer0_outputs(2865));
    layer1_outputs(8474) <= not(layer0_outputs(4984));
    layer1_outputs(8475) <= not(layer0_outputs(4985));
    layer1_outputs(8476) <= (layer0_outputs(1287)) or (layer0_outputs(8299));
    layer1_outputs(8477) <= (layer0_outputs(8918)) or (layer0_outputs(3273));
    layer1_outputs(8478) <= layer0_outputs(7388);
    layer1_outputs(8479) <= not(layer0_outputs(5217)) or (layer0_outputs(5517));
    layer1_outputs(8480) <= not(layer0_outputs(1797));
    layer1_outputs(8481) <= not(layer0_outputs(9176));
    layer1_outputs(8482) <= not(layer0_outputs(9279)) or (layer0_outputs(7125));
    layer1_outputs(8483) <= '0';
    layer1_outputs(8484) <= not(layer0_outputs(1008));
    layer1_outputs(8485) <= not((layer0_outputs(4674)) and (layer0_outputs(8472)));
    layer1_outputs(8486) <= (layer0_outputs(4650)) and not (layer0_outputs(2837));
    layer1_outputs(8487) <= not(layer0_outputs(9025));
    layer1_outputs(8488) <= '0';
    layer1_outputs(8489) <= not(layer0_outputs(4514)) or (layer0_outputs(8206));
    layer1_outputs(8490) <= (layer0_outputs(8686)) and not (layer0_outputs(802));
    layer1_outputs(8491) <= (layer0_outputs(9241)) xor (layer0_outputs(1757));
    layer1_outputs(8492) <= not(layer0_outputs(9635));
    layer1_outputs(8493) <= (layer0_outputs(760)) and not (layer0_outputs(4464));
    layer1_outputs(8494) <= not((layer0_outputs(3339)) or (layer0_outputs(675)));
    layer1_outputs(8495) <= not(layer0_outputs(1331));
    layer1_outputs(8496) <= (layer0_outputs(323)) and (layer0_outputs(1822));
    layer1_outputs(8497) <= not((layer0_outputs(3716)) and (layer0_outputs(5866)));
    layer1_outputs(8498) <= not(layer0_outputs(2547)) or (layer0_outputs(9093));
    layer1_outputs(8499) <= not((layer0_outputs(2898)) and (layer0_outputs(3340)));
    layer1_outputs(8500) <= layer0_outputs(7133);
    layer1_outputs(8501) <= not((layer0_outputs(4852)) and (layer0_outputs(2552)));
    layer1_outputs(8502) <= layer0_outputs(1804);
    layer1_outputs(8503) <= layer0_outputs(6273);
    layer1_outputs(8504) <= not(layer0_outputs(4024));
    layer1_outputs(8505) <= not((layer0_outputs(7167)) and (layer0_outputs(2872)));
    layer1_outputs(8506) <= layer0_outputs(7632);
    layer1_outputs(8507) <= not(layer0_outputs(5276));
    layer1_outputs(8508) <= layer0_outputs(9643);
    layer1_outputs(8509) <= not((layer0_outputs(8386)) and (layer0_outputs(4708)));
    layer1_outputs(8510) <= not((layer0_outputs(181)) or (layer0_outputs(8422)));
    layer1_outputs(8511) <= layer0_outputs(9894);
    layer1_outputs(8512) <= (layer0_outputs(7326)) or (layer0_outputs(3123));
    layer1_outputs(8513) <= '1';
    layer1_outputs(8514) <= layer0_outputs(6998);
    layer1_outputs(8515) <= not(layer0_outputs(9986));
    layer1_outputs(8516) <= layer0_outputs(3537);
    layer1_outputs(8517) <= not(layer0_outputs(4320)) or (layer0_outputs(6456));
    layer1_outputs(8518) <= layer0_outputs(1605);
    layer1_outputs(8519) <= not(layer0_outputs(5906));
    layer1_outputs(8520) <= (layer0_outputs(10064)) xor (layer0_outputs(524));
    layer1_outputs(8521) <= (layer0_outputs(3070)) and not (layer0_outputs(9387));
    layer1_outputs(8522) <= '0';
    layer1_outputs(8523) <= layer0_outputs(7017);
    layer1_outputs(8524) <= layer0_outputs(890);
    layer1_outputs(8525) <= layer0_outputs(1674);
    layer1_outputs(8526) <= not(layer0_outputs(6692)) or (layer0_outputs(2989));
    layer1_outputs(8527) <= not(layer0_outputs(5218));
    layer1_outputs(8528) <= not(layer0_outputs(8399));
    layer1_outputs(8529) <= not(layer0_outputs(3189)) or (layer0_outputs(6108));
    layer1_outputs(8530) <= not(layer0_outputs(6580));
    layer1_outputs(8531) <= (layer0_outputs(1001)) and not (layer0_outputs(439));
    layer1_outputs(8532) <= not((layer0_outputs(4488)) and (layer0_outputs(9644)));
    layer1_outputs(8533) <= not(layer0_outputs(5360)) or (layer0_outputs(8401));
    layer1_outputs(8534) <= layer0_outputs(5452);
    layer1_outputs(8535) <= (layer0_outputs(2178)) or (layer0_outputs(3550));
    layer1_outputs(8536) <= layer0_outputs(2448);
    layer1_outputs(8537) <= (layer0_outputs(3564)) or (layer0_outputs(4758));
    layer1_outputs(8538) <= not((layer0_outputs(2017)) or (layer0_outputs(5475)));
    layer1_outputs(8539) <= (layer0_outputs(6761)) and not (layer0_outputs(7562));
    layer1_outputs(8540) <= (layer0_outputs(1003)) and not (layer0_outputs(9236));
    layer1_outputs(8541) <= layer0_outputs(7934);
    layer1_outputs(8542) <= (layer0_outputs(8142)) or (layer0_outputs(1202));
    layer1_outputs(8543) <= (layer0_outputs(720)) or (layer0_outputs(1327));
    layer1_outputs(8544) <= not(layer0_outputs(6542)) or (layer0_outputs(9461));
    layer1_outputs(8545) <= layer0_outputs(3259);
    layer1_outputs(8546) <= not((layer0_outputs(4588)) or (layer0_outputs(8715)));
    layer1_outputs(8547) <= not(layer0_outputs(7264)) or (layer0_outputs(82));
    layer1_outputs(8548) <= layer0_outputs(321);
    layer1_outputs(8549) <= not((layer0_outputs(986)) and (layer0_outputs(8685)));
    layer1_outputs(8550) <= (layer0_outputs(3361)) and not (layer0_outputs(4638));
    layer1_outputs(8551) <= not((layer0_outputs(3496)) and (layer0_outputs(4848)));
    layer1_outputs(8552) <= layer0_outputs(254);
    layer1_outputs(8553) <= (layer0_outputs(2932)) and not (layer0_outputs(6419));
    layer1_outputs(8554) <= (layer0_outputs(588)) or (layer0_outputs(3797));
    layer1_outputs(8555) <= layer0_outputs(1934);
    layer1_outputs(8556) <= not(layer0_outputs(6231));
    layer1_outputs(8557) <= not((layer0_outputs(7473)) and (layer0_outputs(2523)));
    layer1_outputs(8558) <= not((layer0_outputs(9744)) and (layer0_outputs(1987)));
    layer1_outputs(8559) <= not(layer0_outputs(2226));
    layer1_outputs(8560) <= not((layer0_outputs(5153)) and (layer0_outputs(6192)));
    layer1_outputs(8561) <= not(layer0_outputs(3349)) or (layer0_outputs(1005));
    layer1_outputs(8562) <= not(layer0_outputs(1912)) or (layer0_outputs(4202));
    layer1_outputs(8563) <= not((layer0_outputs(7263)) and (layer0_outputs(2427)));
    layer1_outputs(8564) <= not(layer0_outputs(4757));
    layer1_outputs(8565) <= (layer0_outputs(7555)) and (layer0_outputs(4317));
    layer1_outputs(8566) <= not((layer0_outputs(128)) or (layer0_outputs(1179)));
    layer1_outputs(8567) <= (layer0_outputs(4475)) and not (layer0_outputs(9002));
    layer1_outputs(8568) <= (layer0_outputs(3360)) and not (layer0_outputs(3920));
    layer1_outputs(8569) <= (layer0_outputs(2578)) and not (layer0_outputs(9790));
    layer1_outputs(8570) <= (layer0_outputs(4127)) or (layer0_outputs(8035));
    layer1_outputs(8571) <= not((layer0_outputs(6904)) and (layer0_outputs(833)));
    layer1_outputs(8572) <= not((layer0_outputs(5828)) and (layer0_outputs(1941)));
    layer1_outputs(8573) <= (layer0_outputs(9570)) or (layer0_outputs(4105));
    layer1_outputs(8574) <= (layer0_outputs(1073)) and not (layer0_outputs(8122));
    layer1_outputs(8575) <= not(layer0_outputs(6547)) or (layer0_outputs(8605));
    layer1_outputs(8576) <= layer0_outputs(5000);
    layer1_outputs(8577) <= not(layer0_outputs(2540));
    layer1_outputs(8578) <= not((layer0_outputs(3853)) xor (layer0_outputs(2733)));
    layer1_outputs(8579) <= '0';
    layer1_outputs(8580) <= not(layer0_outputs(4266));
    layer1_outputs(8581) <= (layer0_outputs(7330)) xor (layer0_outputs(845));
    layer1_outputs(8582) <= not(layer0_outputs(9526));
    layer1_outputs(8583) <= (layer0_outputs(2998)) and not (layer0_outputs(6535));
    layer1_outputs(8584) <= (layer0_outputs(1117)) and not (layer0_outputs(9152));
    layer1_outputs(8585) <= (layer0_outputs(8601)) and not (layer0_outputs(5050));
    layer1_outputs(8586) <= (layer0_outputs(5932)) and (layer0_outputs(3271));
    layer1_outputs(8587) <= not(layer0_outputs(5920));
    layer1_outputs(8588) <= '0';
    layer1_outputs(8589) <= layer0_outputs(3566);
    layer1_outputs(8590) <= '1';
    layer1_outputs(8591) <= not((layer0_outputs(7117)) xor (layer0_outputs(4463)));
    layer1_outputs(8592) <= not(layer0_outputs(4383));
    layer1_outputs(8593) <= layer0_outputs(2902);
    layer1_outputs(8594) <= not((layer0_outputs(2489)) or (layer0_outputs(4057)));
    layer1_outputs(8595) <= (layer0_outputs(2780)) xor (layer0_outputs(8098));
    layer1_outputs(8596) <= (layer0_outputs(1299)) and not (layer0_outputs(1392));
    layer1_outputs(8597) <= not(layer0_outputs(5575));
    layer1_outputs(8598) <= (layer0_outputs(4459)) and not (layer0_outputs(4053));
    layer1_outputs(8599) <= not(layer0_outputs(8871)) or (layer0_outputs(3366));
    layer1_outputs(8600) <= not(layer0_outputs(9248)) or (layer0_outputs(6608));
    layer1_outputs(8601) <= (layer0_outputs(3384)) or (layer0_outputs(5560));
    layer1_outputs(8602) <= not(layer0_outputs(7967));
    layer1_outputs(8603) <= not((layer0_outputs(9651)) xor (layer0_outputs(406)));
    layer1_outputs(8604) <= layer0_outputs(7701);
    layer1_outputs(8605) <= '0';
    layer1_outputs(8606) <= (layer0_outputs(9459)) or (layer0_outputs(4105));
    layer1_outputs(8607) <= layer0_outputs(3998);
    layer1_outputs(8608) <= not(layer0_outputs(3552));
    layer1_outputs(8609) <= layer0_outputs(3415);
    layer1_outputs(8610) <= not(layer0_outputs(582)) or (layer0_outputs(1676));
    layer1_outputs(8611) <= (layer0_outputs(4368)) or (layer0_outputs(10015));
    layer1_outputs(8612) <= layer0_outputs(9992);
    layer1_outputs(8613) <= '0';
    layer1_outputs(8614) <= not((layer0_outputs(4304)) or (layer0_outputs(4527)));
    layer1_outputs(8615) <= not((layer0_outputs(5320)) xor (layer0_outputs(2462)));
    layer1_outputs(8616) <= not(layer0_outputs(4365));
    layer1_outputs(8617) <= not((layer0_outputs(245)) and (layer0_outputs(10220)));
    layer1_outputs(8618) <= (layer0_outputs(6948)) and not (layer0_outputs(8448));
    layer1_outputs(8619) <= not(layer0_outputs(352)) or (layer0_outputs(2059));
    layer1_outputs(8620) <= not(layer0_outputs(602));
    layer1_outputs(8621) <= not(layer0_outputs(5921)) or (layer0_outputs(4312));
    layer1_outputs(8622) <= (layer0_outputs(9080)) or (layer0_outputs(4538));
    layer1_outputs(8623) <= not((layer0_outputs(4916)) or (layer0_outputs(9614)));
    layer1_outputs(8624) <= not(layer0_outputs(5284)) or (layer0_outputs(6239));
    layer1_outputs(8625) <= not(layer0_outputs(4431));
    layer1_outputs(8626) <= (layer0_outputs(2201)) or (layer0_outputs(6128));
    layer1_outputs(8627) <= layer0_outputs(681);
    layer1_outputs(8628) <= layer0_outputs(8653);
    layer1_outputs(8629) <= (layer0_outputs(9375)) and not (layer0_outputs(7684));
    layer1_outputs(8630) <= layer0_outputs(9338);
    layer1_outputs(8631) <= not(layer0_outputs(70));
    layer1_outputs(8632) <= not((layer0_outputs(2165)) xor (layer0_outputs(8167)));
    layer1_outputs(8633) <= not(layer0_outputs(917)) or (layer0_outputs(8045));
    layer1_outputs(8634) <= not(layer0_outputs(7201)) or (layer0_outputs(7845));
    layer1_outputs(8635) <= '0';
    layer1_outputs(8636) <= (layer0_outputs(220)) and not (layer0_outputs(6452));
    layer1_outputs(8637) <= not(layer0_outputs(7823)) or (layer0_outputs(6044));
    layer1_outputs(8638) <= (layer0_outputs(7789)) or (layer0_outputs(8998));
    layer1_outputs(8639) <= (layer0_outputs(205)) and not (layer0_outputs(6532));
    layer1_outputs(8640) <= not((layer0_outputs(6367)) or (layer0_outputs(7509)));
    layer1_outputs(8641) <= not(layer0_outputs(4556));
    layer1_outputs(8642) <= not((layer0_outputs(3518)) xor (layer0_outputs(1389)));
    layer1_outputs(8643) <= not(layer0_outputs(4884));
    layer1_outputs(8644) <= not((layer0_outputs(2910)) and (layer0_outputs(3408)));
    layer1_outputs(8645) <= not(layer0_outputs(9315));
    layer1_outputs(8646) <= not(layer0_outputs(2051)) or (layer0_outputs(5570));
    layer1_outputs(8647) <= (layer0_outputs(6080)) xor (layer0_outputs(311));
    layer1_outputs(8648) <= (layer0_outputs(5584)) xor (layer0_outputs(2962));
    layer1_outputs(8649) <= layer0_outputs(7417);
    layer1_outputs(8650) <= '1';
    layer1_outputs(8651) <= layer0_outputs(1482);
    layer1_outputs(8652) <= (layer0_outputs(4995)) xor (layer0_outputs(1926));
    layer1_outputs(8653) <= (layer0_outputs(6742)) and (layer0_outputs(8477));
    layer1_outputs(8654) <= not(layer0_outputs(1037));
    layer1_outputs(8655) <= '1';
    layer1_outputs(8656) <= layer0_outputs(3095);
    layer1_outputs(8657) <= not(layer0_outputs(9650)) or (layer0_outputs(7559));
    layer1_outputs(8658) <= (layer0_outputs(2591)) and (layer0_outputs(2471));
    layer1_outputs(8659) <= not(layer0_outputs(1338));
    layer1_outputs(8660) <= not(layer0_outputs(7122)) or (layer0_outputs(4285));
    layer1_outputs(8661) <= layer0_outputs(1415);
    layer1_outputs(8662) <= not(layer0_outputs(3227));
    layer1_outputs(8663) <= not(layer0_outputs(4908));
    layer1_outputs(8664) <= (layer0_outputs(1175)) or (layer0_outputs(3984));
    layer1_outputs(8665) <= not(layer0_outputs(3949));
    layer1_outputs(8666) <= (layer0_outputs(7475)) xor (layer0_outputs(6185));
    layer1_outputs(8667) <= not(layer0_outputs(768));
    layer1_outputs(8668) <= layer0_outputs(9220);
    layer1_outputs(8669) <= not((layer0_outputs(3835)) or (layer0_outputs(7190)));
    layer1_outputs(8670) <= not(layer0_outputs(5944));
    layer1_outputs(8671) <= not(layer0_outputs(3670)) or (layer0_outputs(5260));
    layer1_outputs(8672) <= not(layer0_outputs(3659));
    layer1_outputs(8673) <= (layer0_outputs(3502)) and (layer0_outputs(8723));
    layer1_outputs(8674) <= not(layer0_outputs(8730));
    layer1_outputs(8675) <= not(layer0_outputs(9158));
    layer1_outputs(8676) <= not(layer0_outputs(3273)) or (layer0_outputs(4933));
    layer1_outputs(8677) <= (layer0_outputs(2605)) and not (layer0_outputs(918));
    layer1_outputs(8678) <= layer0_outputs(2280);
    layer1_outputs(8679) <= not(layer0_outputs(1704));
    layer1_outputs(8680) <= not(layer0_outputs(1742));
    layer1_outputs(8681) <= not(layer0_outputs(1567));
    layer1_outputs(8682) <= not(layer0_outputs(10096));
    layer1_outputs(8683) <= (layer0_outputs(2415)) or (layer0_outputs(1992));
    layer1_outputs(8684) <= layer0_outputs(2946);
    layer1_outputs(8685) <= (layer0_outputs(6910)) or (layer0_outputs(8218));
    layer1_outputs(8686) <= not((layer0_outputs(4128)) or (layer0_outputs(9213)));
    layer1_outputs(8687) <= (layer0_outputs(6327)) and (layer0_outputs(7269));
    layer1_outputs(8688) <= not((layer0_outputs(4925)) or (layer0_outputs(9722)));
    layer1_outputs(8689) <= not((layer0_outputs(4190)) or (layer0_outputs(2097)));
    layer1_outputs(8690) <= not((layer0_outputs(3050)) or (layer0_outputs(2931)));
    layer1_outputs(8691) <= (layer0_outputs(4685)) and not (layer0_outputs(6455));
    layer1_outputs(8692) <= layer0_outputs(7423);
    layer1_outputs(8693) <= layer0_outputs(5193);
    layer1_outputs(8694) <= (layer0_outputs(5729)) and not (layer0_outputs(7583));
    layer1_outputs(8695) <= (layer0_outputs(1644)) and (layer0_outputs(8332));
    layer1_outputs(8696) <= '0';
    layer1_outputs(8697) <= not(layer0_outputs(5729)) or (layer0_outputs(5587));
    layer1_outputs(8698) <= not(layer0_outputs(1523));
    layer1_outputs(8699) <= (layer0_outputs(4607)) and not (layer0_outputs(653));
    layer1_outputs(8700) <= (layer0_outputs(4487)) and not (layer0_outputs(6488));
    layer1_outputs(8701) <= (layer0_outputs(3746)) and (layer0_outputs(5699));
    layer1_outputs(8702) <= layer0_outputs(8404);
    layer1_outputs(8703) <= layer0_outputs(377);
    layer1_outputs(8704) <= layer0_outputs(6936);
    layer1_outputs(8705) <= layer0_outputs(1497);
    layer1_outputs(8706) <= (layer0_outputs(3529)) or (layer0_outputs(5617));
    layer1_outputs(8707) <= not(layer0_outputs(4002));
    layer1_outputs(8708) <= (layer0_outputs(3998)) and not (layer0_outputs(3933));
    layer1_outputs(8709) <= not(layer0_outputs(2965));
    layer1_outputs(8710) <= not(layer0_outputs(513));
    layer1_outputs(8711) <= layer0_outputs(6547);
    layer1_outputs(8712) <= not((layer0_outputs(2205)) and (layer0_outputs(3583)));
    layer1_outputs(8713) <= (layer0_outputs(815)) and (layer0_outputs(3768));
    layer1_outputs(8714) <= '1';
    layer1_outputs(8715) <= (layer0_outputs(7954)) and (layer0_outputs(9656));
    layer1_outputs(8716) <= '1';
    layer1_outputs(8717) <= (layer0_outputs(4168)) or (layer0_outputs(5091));
    layer1_outputs(8718) <= (layer0_outputs(4733)) and not (layer0_outputs(9066));
    layer1_outputs(8719) <= not(layer0_outputs(696));
    layer1_outputs(8720) <= (layer0_outputs(6692)) or (layer0_outputs(7360));
    layer1_outputs(8721) <= not(layer0_outputs(5557));
    layer1_outputs(8722) <= not((layer0_outputs(2084)) or (layer0_outputs(6750)));
    layer1_outputs(8723) <= (layer0_outputs(9554)) and not (layer0_outputs(9098));
    layer1_outputs(8724) <= layer0_outputs(232);
    layer1_outputs(8725) <= layer0_outputs(2166);
    layer1_outputs(8726) <= layer0_outputs(3090);
    layer1_outputs(8727) <= (layer0_outputs(3993)) or (layer0_outputs(8537));
    layer1_outputs(8728) <= not(layer0_outputs(105)) or (layer0_outputs(2301));
    layer1_outputs(8729) <= not(layer0_outputs(8126));
    layer1_outputs(8730) <= (layer0_outputs(4008)) xor (layer0_outputs(9991));
    layer1_outputs(8731) <= not(layer0_outputs(991));
    layer1_outputs(8732) <= not(layer0_outputs(1586)) or (layer0_outputs(9426));
    layer1_outputs(8733) <= layer0_outputs(10110);
    layer1_outputs(8734) <= layer0_outputs(9697);
    layer1_outputs(8735) <= not(layer0_outputs(4001));
    layer1_outputs(8736) <= layer0_outputs(1385);
    layer1_outputs(8737) <= not(layer0_outputs(6764));
    layer1_outputs(8738) <= (layer0_outputs(1672)) and (layer0_outputs(5020));
    layer1_outputs(8739) <= not((layer0_outputs(4569)) or (layer0_outputs(972)));
    layer1_outputs(8740) <= (layer0_outputs(3151)) and (layer0_outputs(8006));
    layer1_outputs(8741) <= layer0_outputs(8572);
    layer1_outputs(8742) <= not(layer0_outputs(8307));
    layer1_outputs(8743) <= (layer0_outputs(1849)) or (layer0_outputs(3985));
    layer1_outputs(8744) <= layer0_outputs(899);
    layer1_outputs(8745) <= (layer0_outputs(6363)) and not (layer0_outputs(4203));
    layer1_outputs(8746) <= (layer0_outputs(8262)) and not (layer0_outputs(6870));
    layer1_outputs(8747) <= not(layer0_outputs(8364)) or (layer0_outputs(7295));
    layer1_outputs(8748) <= not((layer0_outputs(1701)) or (layer0_outputs(9043)));
    layer1_outputs(8749) <= (layer0_outputs(7942)) or (layer0_outputs(296));
    layer1_outputs(8750) <= '1';
    layer1_outputs(8751) <= layer0_outputs(2475);
    layer1_outputs(8752) <= not(layer0_outputs(2907)) or (layer0_outputs(4497));
    layer1_outputs(8753) <= not(layer0_outputs(8290)) or (layer0_outputs(3557));
    layer1_outputs(8754) <= (layer0_outputs(6192)) xor (layer0_outputs(7095));
    layer1_outputs(8755) <= not((layer0_outputs(7521)) or (layer0_outputs(3983)));
    layer1_outputs(8756) <= not(layer0_outputs(9769));
    layer1_outputs(8757) <= not((layer0_outputs(319)) and (layer0_outputs(3866)));
    layer1_outputs(8758) <= not((layer0_outputs(5529)) and (layer0_outputs(9965)));
    layer1_outputs(8759) <= not(layer0_outputs(8603));
    layer1_outputs(8760) <= not(layer0_outputs(7603));
    layer1_outputs(8761) <= not(layer0_outputs(10183)) or (layer0_outputs(1334));
    layer1_outputs(8762) <= not(layer0_outputs(6236));
    layer1_outputs(8763) <= not(layer0_outputs(1028));
    layer1_outputs(8764) <= (layer0_outputs(425)) and (layer0_outputs(1211));
    layer1_outputs(8765) <= not(layer0_outputs(8136));
    layer1_outputs(8766) <= layer0_outputs(5847);
    layer1_outputs(8767) <= not((layer0_outputs(9042)) or (layer0_outputs(3950)));
    layer1_outputs(8768) <= not((layer0_outputs(5824)) and (layer0_outputs(9898)));
    layer1_outputs(8769) <= not(layer0_outputs(1324));
    layer1_outputs(8770) <= not(layer0_outputs(365));
    layer1_outputs(8771) <= layer0_outputs(1372);
    layer1_outputs(8772) <= layer0_outputs(1123);
    layer1_outputs(8773) <= not(layer0_outputs(2739));
    layer1_outputs(8774) <= not(layer0_outputs(59));
    layer1_outputs(8775) <= not((layer0_outputs(9836)) xor (layer0_outputs(3324)));
    layer1_outputs(8776) <= layer0_outputs(6673);
    layer1_outputs(8777) <= layer0_outputs(1984);
    layer1_outputs(8778) <= (layer0_outputs(5543)) and not (layer0_outputs(1486));
    layer1_outputs(8779) <= not(layer0_outputs(2921));
    layer1_outputs(8780) <= not(layer0_outputs(296));
    layer1_outputs(8781) <= (layer0_outputs(2255)) xor (layer0_outputs(4838));
    layer1_outputs(8782) <= layer0_outputs(5382);
    layer1_outputs(8783) <= (layer0_outputs(3913)) and not (layer0_outputs(5952));
    layer1_outputs(8784) <= not(layer0_outputs(148));
    layer1_outputs(8785) <= not(layer0_outputs(9182));
    layer1_outputs(8786) <= not(layer0_outputs(4504)) or (layer0_outputs(1142));
    layer1_outputs(8787) <= (layer0_outputs(3694)) and (layer0_outputs(9656));
    layer1_outputs(8788) <= '1';
    layer1_outputs(8789) <= not((layer0_outputs(831)) or (layer0_outputs(8610)));
    layer1_outputs(8790) <= layer0_outputs(6951);
    layer1_outputs(8791) <= layer0_outputs(340);
    layer1_outputs(8792) <= (layer0_outputs(9948)) and not (layer0_outputs(1978));
    layer1_outputs(8793) <= not(layer0_outputs(5469)) or (layer0_outputs(636));
    layer1_outputs(8794) <= not((layer0_outputs(1010)) and (layer0_outputs(3327)));
    layer1_outputs(8795) <= layer0_outputs(9356);
    layer1_outputs(8796) <= not(layer0_outputs(5194));
    layer1_outputs(8797) <= not(layer0_outputs(4134));
    layer1_outputs(8798) <= (layer0_outputs(72)) and not (layer0_outputs(260));
    layer1_outputs(8799) <= layer0_outputs(1896);
    layer1_outputs(8800) <= not(layer0_outputs(328)) or (layer0_outputs(5153));
    layer1_outputs(8801) <= layer0_outputs(1436);
    layer1_outputs(8802) <= (layer0_outputs(7196)) and not (layer0_outputs(2855));
    layer1_outputs(8803) <= not(layer0_outputs(259));
    layer1_outputs(8804) <= not(layer0_outputs(1134));
    layer1_outputs(8805) <= (layer0_outputs(4723)) xor (layer0_outputs(7483));
    layer1_outputs(8806) <= layer0_outputs(530);
    layer1_outputs(8807) <= layer0_outputs(5138);
    layer1_outputs(8808) <= not(layer0_outputs(182));
    layer1_outputs(8809) <= not((layer0_outputs(4980)) or (layer0_outputs(433)));
    layer1_outputs(8810) <= layer0_outputs(6241);
    layer1_outputs(8811) <= (layer0_outputs(7226)) or (layer0_outputs(2764));
    layer1_outputs(8812) <= (layer0_outputs(3816)) and not (layer0_outputs(5609));
    layer1_outputs(8813) <= (layer0_outputs(6314)) and not (layer0_outputs(979));
    layer1_outputs(8814) <= not(layer0_outputs(9422));
    layer1_outputs(8815) <= not(layer0_outputs(10164));
    layer1_outputs(8816) <= not((layer0_outputs(287)) and (layer0_outputs(1655)));
    layer1_outputs(8817) <= layer0_outputs(8121);
    layer1_outputs(8818) <= not(layer0_outputs(1484));
    layer1_outputs(8819) <= not(layer0_outputs(306)) or (layer0_outputs(3569));
    layer1_outputs(8820) <= (layer0_outputs(4187)) and not (layer0_outputs(6173));
    layer1_outputs(8821) <= layer0_outputs(3390);
    layer1_outputs(8822) <= (layer0_outputs(6890)) xor (layer0_outputs(5930));
    layer1_outputs(8823) <= layer0_outputs(4603);
    layer1_outputs(8824) <= layer0_outputs(4836);
    layer1_outputs(8825) <= not((layer0_outputs(4984)) and (layer0_outputs(3625)));
    layer1_outputs(8826) <= not(layer0_outputs(7542));
    layer1_outputs(8827) <= not((layer0_outputs(6343)) and (layer0_outputs(8146)));
    layer1_outputs(8828) <= (layer0_outputs(9257)) and not (layer0_outputs(9592));
    layer1_outputs(8829) <= not(layer0_outputs(4501)) or (layer0_outputs(1520));
    layer1_outputs(8830) <= (layer0_outputs(6748)) and not (layer0_outputs(1664));
    layer1_outputs(8831) <= (layer0_outputs(7414)) xor (layer0_outputs(8495));
    layer1_outputs(8832) <= not((layer0_outputs(168)) and (layer0_outputs(1638)));
    layer1_outputs(8833) <= (layer0_outputs(3493)) and not (layer0_outputs(9266));
    layer1_outputs(8834) <= layer0_outputs(692);
    layer1_outputs(8835) <= '1';
    layer1_outputs(8836) <= '1';
    layer1_outputs(8837) <= not(layer0_outputs(1929));
    layer1_outputs(8838) <= (layer0_outputs(9107)) and not (layer0_outputs(1303));
    layer1_outputs(8839) <= layer0_outputs(6234);
    layer1_outputs(8840) <= (layer0_outputs(8324)) or (layer0_outputs(4947));
    layer1_outputs(8841) <= layer0_outputs(1320);
    layer1_outputs(8842) <= (layer0_outputs(5619)) and not (layer0_outputs(8733));
    layer1_outputs(8843) <= not(layer0_outputs(8578)) or (layer0_outputs(818));
    layer1_outputs(8844) <= not((layer0_outputs(9707)) and (layer0_outputs(10189)));
    layer1_outputs(8845) <= (layer0_outputs(6165)) and not (layer0_outputs(5130));
    layer1_outputs(8846) <= not(layer0_outputs(155));
    layer1_outputs(8847) <= layer0_outputs(9907);
    layer1_outputs(8848) <= not(layer0_outputs(225));
    layer1_outputs(8849) <= '1';
    layer1_outputs(8850) <= layer0_outputs(9924);
    layer1_outputs(8851) <= layer0_outputs(7312);
    layer1_outputs(8852) <= not(layer0_outputs(821));
    layer1_outputs(8853) <= (layer0_outputs(7211)) and (layer0_outputs(4874));
    layer1_outputs(8854) <= not(layer0_outputs(1799)) or (layer0_outputs(2718));
    layer1_outputs(8855) <= not((layer0_outputs(1629)) and (layer0_outputs(7261)));
    layer1_outputs(8856) <= not(layer0_outputs(7593));
    layer1_outputs(8857) <= layer0_outputs(9703);
    layer1_outputs(8858) <= not((layer0_outputs(3130)) or (layer0_outputs(3300)));
    layer1_outputs(8859) <= not(layer0_outputs(612)) or (layer0_outputs(2311));
    layer1_outputs(8860) <= not(layer0_outputs(202));
    layer1_outputs(8861) <= not(layer0_outputs(7868));
    layer1_outputs(8862) <= not((layer0_outputs(4119)) and (layer0_outputs(7380)));
    layer1_outputs(8863) <= layer0_outputs(8468);
    layer1_outputs(8864) <= layer0_outputs(9324);
    layer1_outputs(8865) <= (layer0_outputs(2463)) and not (layer0_outputs(2329));
    layer1_outputs(8866) <= (layer0_outputs(9100)) or (layer0_outputs(10074));
    layer1_outputs(8867) <= layer0_outputs(8336);
    layer1_outputs(8868) <= not((layer0_outputs(8984)) and (layer0_outputs(4307)));
    layer1_outputs(8869) <= not((layer0_outputs(2408)) and (layer0_outputs(4340)));
    layer1_outputs(8870) <= not(layer0_outputs(8207));
    layer1_outputs(8871) <= '0';
    layer1_outputs(8872) <= not(layer0_outputs(7153)) or (layer0_outputs(4382));
    layer1_outputs(8873) <= layer0_outputs(1013);
    layer1_outputs(8874) <= (layer0_outputs(8904)) xor (layer0_outputs(9978));
    layer1_outputs(8875) <= (layer0_outputs(4508)) and (layer0_outputs(10203));
    layer1_outputs(8876) <= not(layer0_outputs(2539)) or (layer0_outputs(2048));
    layer1_outputs(8877) <= not(layer0_outputs(1749));
    layer1_outputs(8878) <= (layer0_outputs(8298)) and not (layer0_outputs(186));
    layer1_outputs(8879) <= not((layer0_outputs(6822)) and (layer0_outputs(2551)));
    layer1_outputs(8880) <= not((layer0_outputs(3091)) or (layer0_outputs(10153)));
    layer1_outputs(8881) <= layer0_outputs(3449);
    layer1_outputs(8882) <= layer0_outputs(5711);
    layer1_outputs(8883) <= not(layer0_outputs(5624));
    layer1_outputs(8884) <= not((layer0_outputs(7916)) and (layer0_outputs(3179)));
    layer1_outputs(8885) <= not((layer0_outputs(4615)) or (layer0_outputs(3979)));
    layer1_outputs(8886) <= not(layer0_outputs(2114));
    layer1_outputs(8887) <= (layer0_outputs(7265)) and not (layer0_outputs(5157));
    layer1_outputs(8888) <= (layer0_outputs(7833)) and not (layer0_outputs(9405));
    layer1_outputs(8889) <= layer0_outputs(2273);
    layer1_outputs(8890) <= (layer0_outputs(9918)) and not (layer0_outputs(6043));
    layer1_outputs(8891) <= layer0_outputs(3563);
    layer1_outputs(8892) <= (layer0_outputs(3662)) or (layer0_outputs(7903));
    layer1_outputs(8893) <= (layer0_outputs(2609)) and not (layer0_outputs(2854));
    layer1_outputs(8894) <= (layer0_outputs(681)) xor (layer0_outputs(2591));
    layer1_outputs(8895) <= not(layer0_outputs(6701)) or (layer0_outputs(10033));
    layer1_outputs(8896) <= not(layer0_outputs(7141));
    layer1_outputs(8897) <= (layer0_outputs(2853)) and (layer0_outputs(1168));
    layer1_outputs(8898) <= (layer0_outputs(6265)) and not (layer0_outputs(1942));
    layer1_outputs(8899) <= not(layer0_outputs(8977)) or (layer0_outputs(4372));
    layer1_outputs(8900) <= not(layer0_outputs(9623)) or (layer0_outputs(4778));
    layer1_outputs(8901) <= layer0_outputs(6084);
    layer1_outputs(8902) <= (layer0_outputs(427)) and not (layer0_outputs(3331));
    layer1_outputs(8903) <= not(layer0_outputs(5068)) or (layer0_outputs(3818));
    layer1_outputs(8904) <= (layer0_outputs(4298)) or (layer0_outputs(4701));
    layer1_outputs(8905) <= (layer0_outputs(3463)) or (layer0_outputs(9709));
    layer1_outputs(8906) <= not(layer0_outputs(5826)) or (layer0_outputs(4090));
    layer1_outputs(8907) <= layer0_outputs(6421);
    layer1_outputs(8908) <= not(layer0_outputs(3517)) or (layer0_outputs(4084));
    layer1_outputs(8909) <= not(layer0_outputs(4027));
    layer1_outputs(8910) <= (layer0_outputs(4854)) xor (layer0_outputs(8345));
    layer1_outputs(8911) <= (layer0_outputs(6147)) xor (layer0_outputs(6989));
    layer1_outputs(8912) <= not((layer0_outputs(6742)) and (layer0_outputs(8429)));
    layer1_outputs(8913) <= layer0_outputs(12);
    layer1_outputs(8914) <= (layer0_outputs(6114)) and not (layer0_outputs(8057));
    layer1_outputs(8915) <= not((layer0_outputs(7374)) xor (layer0_outputs(7964)));
    layer1_outputs(8916) <= (layer0_outputs(298)) and (layer0_outputs(2523));
    layer1_outputs(8917) <= not(layer0_outputs(4450)) or (layer0_outputs(10207));
    layer1_outputs(8918) <= layer0_outputs(6874);
    layer1_outputs(8919) <= not((layer0_outputs(8371)) or (layer0_outputs(5296)));
    layer1_outputs(8920) <= not((layer0_outputs(6212)) or (layer0_outputs(8512)));
    layer1_outputs(8921) <= layer0_outputs(5383);
    layer1_outputs(8922) <= not(layer0_outputs(2704)) or (layer0_outputs(10141));
    layer1_outputs(8923) <= (layer0_outputs(6839)) xor (layer0_outputs(2003));
    layer1_outputs(8924) <= not((layer0_outputs(2786)) or (layer0_outputs(3381)));
    layer1_outputs(8925) <= not(layer0_outputs(5559));
    layer1_outputs(8926) <= layer0_outputs(1631);
    layer1_outputs(8927) <= (layer0_outputs(6678)) or (layer0_outputs(1138));
    layer1_outputs(8928) <= (layer0_outputs(7110)) xor (layer0_outputs(3853));
    layer1_outputs(8929) <= not((layer0_outputs(3477)) and (layer0_outputs(8693)));
    layer1_outputs(8930) <= layer0_outputs(3898);
    layer1_outputs(8931) <= not((layer0_outputs(1977)) and (layer0_outputs(4903)));
    layer1_outputs(8932) <= layer0_outputs(4764);
    layer1_outputs(8933) <= layer0_outputs(4373);
    layer1_outputs(8934) <= (layer0_outputs(4358)) or (layer0_outputs(1501));
    layer1_outputs(8935) <= not((layer0_outputs(3533)) xor (layer0_outputs(6403)));
    layer1_outputs(8936) <= not(layer0_outputs(2939));
    layer1_outputs(8937) <= (layer0_outputs(2656)) and not (layer0_outputs(462));
    layer1_outputs(8938) <= layer0_outputs(1960);
    layer1_outputs(8939) <= (layer0_outputs(9495)) xor (layer0_outputs(7538));
    layer1_outputs(8940) <= not((layer0_outputs(4745)) and (layer0_outputs(5520)));
    layer1_outputs(8941) <= not(layer0_outputs(6100)) or (layer0_outputs(3917));
    layer1_outputs(8942) <= (layer0_outputs(2868)) and not (layer0_outputs(6035));
    layer1_outputs(8943) <= (layer0_outputs(3551)) or (layer0_outputs(6163));
    layer1_outputs(8944) <= not((layer0_outputs(1454)) or (layer0_outputs(4592)));
    layer1_outputs(8945) <= not(layer0_outputs(1666)) or (layer0_outputs(8076));
    layer1_outputs(8946) <= not(layer0_outputs(6905));
    layer1_outputs(8947) <= not(layer0_outputs(2537));
    layer1_outputs(8948) <= not((layer0_outputs(1566)) and (layer0_outputs(8421)));
    layer1_outputs(8949) <= not((layer0_outputs(3925)) xor (layer0_outputs(690)));
    layer1_outputs(8950) <= not((layer0_outputs(6546)) xor (layer0_outputs(8745)));
    layer1_outputs(8951) <= (layer0_outputs(9812)) and not (layer0_outputs(9135));
    layer1_outputs(8952) <= not(layer0_outputs(8104));
    layer1_outputs(8953) <= layer0_outputs(5951);
    layer1_outputs(8954) <= (layer0_outputs(7017)) and not (layer0_outputs(6171));
    layer1_outputs(8955) <= layer0_outputs(7081);
    layer1_outputs(8956) <= layer0_outputs(2579);
    layer1_outputs(8957) <= not(layer0_outputs(3915));
    layer1_outputs(8958) <= layer0_outputs(6158);
    layer1_outputs(8959) <= not(layer0_outputs(60));
    layer1_outputs(8960) <= not((layer0_outputs(3800)) and (layer0_outputs(9769)));
    layer1_outputs(8961) <= (layer0_outputs(8293)) and (layer0_outputs(5475));
    layer1_outputs(8962) <= layer0_outputs(8373);
    layer1_outputs(8963) <= not(layer0_outputs(6946)) or (layer0_outputs(4057));
    layer1_outputs(8964) <= not((layer0_outputs(2875)) or (layer0_outputs(5356)));
    layer1_outputs(8965) <= not(layer0_outputs(2627));
    layer1_outputs(8966) <= not(layer0_outputs(6381));
    layer1_outputs(8967) <= (layer0_outputs(8771)) and not (layer0_outputs(6644));
    layer1_outputs(8968) <= (layer0_outputs(8730)) or (layer0_outputs(9708));
    layer1_outputs(8969) <= layer0_outputs(9540);
    layer1_outputs(8970) <= layer0_outputs(4406);
    layer1_outputs(8971) <= not(layer0_outputs(5330));
    layer1_outputs(8972) <= not(layer0_outputs(883)) or (layer0_outputs(7793));
    layer1_outputs(8973) <= layer0_outputs(522);
    layer1_outputs(8974) <= layer0_outputs(8169);
    layer1_outputs(8975) <= not(layer0_outputs(2968));
    layer1_outputs(8976) <= not(layer0_outputs(9915));
    layer1_outputs(8977) <= (layer0_outputs(984)) and (layer0_outputs(9745));
    layer1_outputs(8978) <= not(layer0_outputs(6860)) or (layer0_outputs(4647));
    layer1_outputs(8979) <= layer0_outputs(6808);
    layer1_outputs(8980) <= (layer0_outputs(1283)) and not (layer0_outputs(3452));
    layer1_outputs(8981) <= not(layer0_outputs(5230));
    layer1_outputs(8982) <= '1';
    layer1_outputs(8983) <= (layer0_outputs(533)) and not (layer0_outputs(7766));
    layer1_outputs(8984) <= not((layer0_outputs(3287)) and (layer0_outputs(8637)));
    layer1_outputs(8985) <= not(layer0_outputs(4564));
    layer1_outputs(8986) <= (layer0_outputs(8311)) or (layer0_outputs(5169));
    layer1_outputs(8987) <= not(layer0_outputs(4847)) or (layer0_outputs(4399));
    layer1_outputs(8988) <= not((layer0_outputs(1547)) xor (layer0_outputs(5176)));
    layer1_outputs(8989) <= (layer0_outputs(4652)) and (layer0_outputs(4614));
    layer1_outputs(8990) <= (layer0_outputs(3891)) or (layer0_outputs(7271));
    layer1_outputs(8991) <= not(layer0_outputs(5686));
    layer1_outputs(8992) <= not((layer0_outputs(7292)) and (layer0_outputs(6173)));
    layer1_outputs(8993) <= (layer0_outputs(6296)) and not (layer0_outputs(8877));
    layer1_outputs(8994) <= not(layer0_outputs(3654));
    layer1_outputs(8995) <= not(layer0_outputs(2272));
    layer1_outputs(8996) <= not((layer0_outputs(8617)) and (layer0_outputs(9729)));
    layer1_outputs(8997) <= not(layer0_outputs(8096));
    layer1_outputs(8998) <= not(layer0_outputs(7109)) or (layer0_outputs(6260));
    layer1_outputs(8999) <= (layer0_outputs(9813)) xor (layer0_outputs(580));
    layer1_outputs(9000) <= not(layer0_outputs(1151));
    layer1_outputs(9001) <= layer0_outputs(4394);
    layer1_outputs(9002) <= (layer0_outputs(1839)) xor (layer0_outputs(8082));
    layer1_outputs(9003) <= not(layer0_outputs(1841)) or (layer0_outputs(9714));
    layer1_outputs(9004) <= (layer0_outputs(786)) and not (layer0_outputs(1922));
    layer1_outputs(9005) <= (layer0_outputs(7304)) and not (layer0_outputs(8782));
    layer1_outputs(9006) <= layer0_outputs(990);
    layer1_outputs(9007) <= layer0_outputs(8827);
    layer1_outputs(9008) <= not(layer0_outputs(4654));
    layer1_outputs(9009) <= (layer0_outputs(6884)) and not (layer0_outputs(4668));
    layer1_outputs(9010) <= layer0_outputs(8220);
    layer1_outputs(9011) <= (layer0_outputs(7665)) and (layer0_outputs(8600));
    layer1_outputs(9012) <= not(layer0_outputs(5028));
    layer1_outputs(9013) <= (layer0_outputs(3830)) and not (layer0_outputs(478));
    layer1_outputs(9014) <= not(layer0_outputs(7493)) or (layer0_outputs(3008));
    layer1_outputs(9015) <= not(layer0_outputs(8135)) or (layer0_outputs(8755));
    layer1_outputs(9016) <= (layer0_outputs(2016)) and (layer0_outputs(8557));
    layer1_outputs(9017) <= (layer0_outputs(3246)) and not (layer0_outputs(1745));
    layer1_outputs(9018) <= (layer0_outputs(1862)) and (layer0_outputs(6530));
    layer1_outputs(9019) <= '0';
    layer1_outputs(9020) <= not((layer0_outputs(3313)) and (layer0_outputs(449)));
    layer1_outputs(9021) <= not(layer0_outputs(5084));
    layer1_outputs(9022) <= (layer0_outputs(1521)) and not (layer0_outputs(6513));
    layer1_outputs(9023) <= not(layer0_outputs(152));
    layer1_outputs(9024) <= not((layer0_outputs(4385)) and (layer0_outputs(6618)));
    layer1_outputs(9025) <= not(layer0_outputs(10132)) or (layer0_outputs(2326));
    layer1_outputs(9026) <= (layer0_outputs(9984)) or (layer0_outputs(442));
    layer1_outputs(9027) <= (layer0_outputs(5972)) and not (layer0_outputs(9555));
    layer1_outputs(9028) <= not(layer0_outputs(5687));
    layer1_outputs(9029) <= not(layer0_outputs(8567));
    layer1_outputs(9030) <= (layer0_outputs(2844)) and not (layer0_outputs(5509));
    layer1_outputs(9031) <= not(layer0_outputs(7622));
    layer1_outputs(9032) <= not((layer0_outputs(8594)) and (layer0_outputs(9137)));
    layer1_outputs(9033) <= layer0_outputs(7853);
    layer1_outputs(9034) <= not(layer0_outputs(1231));
    layer1_outputs(9035) <= (layer0_outputs(9418)) or (layer0_outputs(6443));
    layer1_outputs(9036) <= (layer0_outputs(8022)) xor (layer0_outputs(9508));
    layer1_outputs(9037) <= not(layer0_outputs(8419));
    layer1_outputs(9038) <= not((layer0_outputs(3113)) or (layer0_outputs(1242)));
    layer1_outputs(9039) <= layer0_outputs(9783);
    layer1_outputs(9040) <= '0';
    layer1_outputs(9041) <= not(layer0_outputs(97));
    layer1_outputs(9042) <= layer0_outputs(9052);
    layer1_outputs(9043) <= layer0_outputs(3092);
    layer1_outputs(9044) <= not(layer0_outputs(9693));
    layer1_outputs(9045) <= not((layer0_outputs(1221)) xor (layer0_outputs(5015)));
    layer1_outputs(9046) <= layer0_outputs(7729);
    layer1_outputs(9047) <= not(layer0_outputs(8023)) or (layer0_outputs(5428));
    layer1_outputs(9048) <= not(layer0_outputs(1751));
    layer1_outputs(9049) <= (layer0_outputs(5656)) and not (layer0_outputs(3080));
    layer1_outputs(9050) <= (layer0_outputs(3348)) and not (layer0_outputs(9627));
    layer1_outputs(9051) <= not((layer0_outputs(9682)) or (layer0_outputs(3009)));
    layer1_outputs(9052) <= (layer0_outputs(2506)) and not (layer0_outputs(2201));
    layer1_outputs(9053) <= not(layer0_outputs(9085));
    layer1_outputs(9054) <= not((layer0_outputs(7470)) and (layer0_outputs(4779)));
    layer1_outputs(9055) <= (layer0_outputs(7460)) xor (layer0_outputs(1458));
    layer1_outputs(9056) <= not((layer0_outputs(5995)) or (layer0_outputs(899)));
    layer1_outputs(9057) <= (layer0_outputs(9789)) and (layer0_outputs(2323));
    layer1_outputs(9058) <= layer0_outputs(1143);
    layer1_outputs(9059) <= layer0_outputs(4413);
    layer1_outputs(9060) <= (layer0_outputs(8461)) and not (layer0_outputs(4706));
    layer1_outputs(9061) <= not((layer0_outputs(2326)) and (layer0_outputs(1652)));
    layer1_outputs(9062) <= (layer0_outputs(6188)) and not (layer0_outputs(3571));
    layer1_outputs(9063) <= not((layer0_outputs(2304)) xor (layer0_outputs(8696)));
    layer1_outputs(9064) <= not(layer0_outputs(76)) or (layer0_outputs(4958));
    layer1_outputs(9065) <= (layer0_outputs(5610)) and (layer0_outputs(4321));
    layer1_outputs(9066) <= (layer0_outputs(972)) or (layer0_outputs(4997));
    layer1_outputs(9067) <= layer0_outputs(10191);
    layer1_outputs(9068) <= not(layer0_outputs(6983));
    layer1_outputs(9069) <= not((layer0_outputs(6583)) or (layer0_outputs(10228)));
    layer1_outputs(9070) <= not(layer0_outputs(1068));
    layer1_outputs(9071) <= not(layer0_outputs(7115));
    layer1_outputs(9072) <= not(layer0_outputs(5753)) or (layer0_outputs(960));
    layer1_outputs(9073) <= (layer0_outputs(8327)) xor (layer0_outputs(574));
    layer1_outputs(9074) <= not(layer0_outputs(6672)) or (layer0_outputs(1160));
    layer1_outputs(9075) <= (layer0_outputs(3065)) or (layer0_outputs(5640));
    layer1_outputs(9076) <= not(layer0_outputs(6338));
    layer1_outputs(9077) <= layer0_outputs(5098);
    layer1_outputs(9078) <= not(layer0_outputs(7586));
    layer1_outputs(9079) <= not(layer0_outputs(9049)) or (layer0_outputs(6868));
    layer1_outputs(9080) <= layer0_outputs(1461);
    layer1_outputs(9081) <= not(layer0_outputs(9916));
    layer1_outputs(9082) <= (layer0_outputs(386)) and (layer0_outputs(9539));
    layer1_outputs(9083) <= not(layer0_outputs(6673)) or (layer0_outputs(1814));
    layer1_outputs(9084) <= layer0_outputs(1201);
    layer1_outputs(9085) <= (layer0_outputs(8412)) xor (layer0_outputs(3709));
    layer1_outputs(9086) <= (layer0_outputs(446)) and not (layer0_outputs(7301));
    layer1_outputs(9087) <= (layer0_outputs(1635)) or (layer0_outputs(8474));
    layer1_outputs(9088) <= layer0_outputs(8263);
    layer1_outputs(9089) <= '1';
    layer1_outputs(9090) <= not(layer0_outputs(2965)) or (layer0_outputs(1761));
    layer1_outputs(9091) <= (layer0_outputs(1684)) or (layer0_outputs(4560));
    layer1_outputs(9092) <= '0';
    layer1_outputs(9093) <= not(layer0_outputs(2033));
    layer1_outputs(9094) <= not((layer0_outputs(3083)) and (layer0_outputs(1598)));
    layer1_outputs(9095) <= layer0_outputs(5764);
    layer1_outputs(9096) <= not(layer0_outputs(10199)) or (layer0_outputs(1286));
    layer1_outputs(9097) <= layer0_outputs(1525);
    layer1_outputs(9098) <= (layer0_outputs(9268)) and not (layer0_outputs(4094));
    layer1_outputs(9099) <= not(layer0_outputs(7541)) or (layer0_outputs(6998));
    layer1_outputs(9100) <= not((layer0_outputs(5050)) xor (layer0_outputs(5086)));
    layer1_outputs(9101) <= not(layer0_outputs(5079)) or (layer0_outputs(3225));
    layer1_outputs(9102) <= not(layer0_outputs(9760));
    layer1_outputs(9103) <= not((layer0_outputs(3402)) or (layer0_outputs(676)));
    layer1_outputs(9104) <= not(layer0_outputs(7448));
    layer1_outputs(9105) <= layer0_outputs(5742);
    layer1_outputs(9106) <= layer0_outputs(3510);
    layer1_outputs(9107) <= (layer0_outputs(6743)) and (layer0_outputs(926));
    layer1_outputs(9108) <= not(layer0_outputs(641));
    layer1_outputs(9109) <= layer0_outputs(7892);
    layer1_outputs(9110) <= (layer0_outputs(9813)) and not (layer0_outputs(5213));
    layer1_outputs(9111) <= '1';
    layer1_outputs(9112) <= (layer0_outputs(6648)) xor (layer0_outputs(4987));
    layer1_outputs(9113) <= (layer0_outputs(5051)) xor (layer0_outputs(7547));
    layer1_outputs(9114) <= layer0_outputs(2682);
    layer1_outputs(9115) <= (layer0_outputs(4855)) xor (layer0_outputs(6985));
    layer1_outputs(9116) <= not((layer0_outputs(2700)) and (layer0_outputs(584)));
    layer1_outputs(9117) <= layer0_outputs(678);
    layer1_outputs(9118) <= not((layer0_outputs(6031)) and (layer0_outputs(8747)));
    layer1_outputs(9119) <= not(layer0_outputs(8036));
    layer1_outputs(9120) <= not((layer0_outputs(7055)) or (layer0_outputs(8562)));
    layer1_outputs(9121) <= not(layer0_outputs(1902)) or (layer0_outputs(8953));
    layer1_outputs(9122) <= not((layer0_outputs(1747)) and (layer0_outputs(538)));
    layer1_outputs(9123) <= not((layer0_outputs(7494)) or (layer0_outputs(8281)));
    layer1_outputs(9124) <= not(layer0_outputs(6925)) or (layer0_outputs(609));
    layer1_outputs(9125) <= (layer0_outputs(468)) and not (layer0_outputs(77));
    layer1_outputs(9126) <= not(layer0_outputs(3912)) or (layer0_outputs(2377));
    layer1_outputs(9127) <= not((layer0_outputs(3595)) or (layer0_outputs(4053)));
    layer1_outputs(9128) <= '0';
    layer1_outputs(9129) <= not((layer0_outputs(10196)) and (layer0_outputs(2389)));
    layer1_outputs(9130) <= (layer0_outputs(6150)) and not (layer0_outputs(6670));
    layer1_outputs(9131) <= layer0_outputs(673);
    layer1_outputs(9132) <= layer0_outputs(2546);
    layer1_outputs(9133) <= (layer0_outputs(8306)) and not (layer0_outputs(4117));
    layer1_outputs(9134) <= not(layer0_outputs(2314));
    layer1_outputs(9135) <= not(layer0_outputs(5550)) or (layer0_outputs(1837));
    layer1_outputs(9136) <= not(layer0_outputs(9423));
    layer1_outputs(9137) <= not((layer0_outputs(653)) xor (layer0_outputs(8695)));
    layer1_outputs(9138) <= layer0_outputs(6902);
    layer1_outputs(9139) <= not(layer0_outputs(7644)) or (layer0_outputs(383));
    layer1_outputs(9140) <= not(layer0_outputs(4601));
    layer1_outputs(9141) <= not(layer0_outputs(1737));
    layer1_outputs(9142) <= (layer0_outputs(2042)) and not (layer0_outputs(7860));
    layer1_outputs(9143) <= '0';
    layer1_outputs(9144) <= layer0_outputs(9445);
    layer1_outputs(9145) <= '1';
    layer1_outputs(9146) <= not(layer0_outputs(8360));
    layer1_outputs(9147) <= (layer0_outputs(2556)) and not (layer0_outputs(6625));
    layer1_outputs(9148) <= (layer0_outputs(3077)) and (layer0_outputs(2661));
    layer1_outputs(9149) <= layer0_outputs(7124);
    layer1_outputs(9150) <= layer0_outputs(2313);
    layer1_outputs(9151) <= not(layer0_outputs(7457)) or (layer0_outputs(3693));
    layer1_outputs(9152) <= (layer0_outputs(987)) and not (layer0_outputs(2500));
    layer1_outputs(9153) <= not(layer0_outputs(7588));
    layer1_outputs(9154) <= not(layer0_outputs(1245));
    layer1_outputs(9155) <= not((layer0_outputs(5548)) xor (layer0_outputs(5568)));
    layer1_outputs(9156) <= (layer0_outputs(7664)) and not (layer0_outputs(6529));
    layer1_outputs(9157) <= (layer0_outputs(2477)) and not (layer0_outputs(4044));
    layer1_outputs(9158) <= layer0_outputs(2650);
    layer1_outputs(9159) <= (layer0_outputs(8923)) xor (layer0_outputs(492));
    layer1_outputs(9160) <= not((layer0_outputs(306)) and (layer0_outputs(5531)));
    layer1_outputs(9161) <= layer0_outputs(3626);
    layer1_outputs(9162) <= layer0_outputs(8073);
    layer1_outputs(9163) <= not(layer0_outputs(6999)) or (layer0_outputs(420));
    layer1_outputs(9164) <= layer0_outputs(3969);
    layer1_outputs(9165) <= (layer0_outputs(7918)) and (layer0_outputs(7368));
    layer1_outputs(9166) <= not((layer0_outputs(7228)) or (layer0_outputs(2651)));
    layer1_outputs(9167) <= (layer0_outputs(1546)) or (layer0_outputs(1718));
    layer1_outputs(9168) <= (layer0_outputs(7605)) and not (layer0_outputs(3455));
    layer1_outputs(9169) <= layer0_outputs(6799);
    layer1_outputs(9170) <= layer0_outputs(2324);
    layer1_outputs(9171) <= layer0_outputs(10224);
    layer1_outputs(9172) <= not(layer0_outputs(6864));
    layer1_outputs(9173) <= not(layer0_outputs(3809));
    layer1_outputs(9174) <= (layer0_outputs(9526)) and (layer0_outputs(764));
    layer1_outputs(9175) <= not(layer0_outputs(2338));
    layer1_outputs(9176) <= layer0_outputs(1528);
    layer1_outputs(9177) <= (layer0_outputs(6757)) xor (layer0_outputs(10046));
    layer1_outputs(9178) <= layer0_outputs(5823);
    layer1_outputs(9179) <= not(layer0_outputs(8558)) or (layer0_outputs(3896));
    layer1_outputs(9180) <= not(layer0_outputs(9928));
    layer1_outputs(9181) <= not(layer0_outputs(3001));
    layer1_outputs(9182) <= not((layer0_outputs(6680)) xor (layer0_outputs(2322)));
    layer1_outputs(9183) <= '0';
    layer1_outputs(9184) <= layer0_outputs(8606);
    layer1_outputs(9185) <= (layer0_outputs(2728)) and not (layer0_outputs(5082));
    layer1_outputs(9186) <= (layer0_outputs(1059)) or (layer0_outputs(2736));
    layer1_outputs(9187) <= not(layer0_outputs(3958));
    layer1_outputs(9188) <= not((layer0_outputs(7989)) and (layer0_outputs(6932)));
    layer1_outputs(9189) <= (layer0_outputs(1808)) xor (layer0_outputs(9139));
    layer1_outputs(9190) <= layer0_outputs(2558);
    layer1_outputs(9191) <= not((layer0_outputs(4138)) xor (layer0_outputs(4961)));
    layer1_outputs(9192) <= (layer0_outputs(5013)) or (layer0_outputs(7927));
    layer1_outputs(9193) <= not(layer0_outputs(9669));
    layer1_outputs(9194) <= not((layer0_outputs(7933)) and (layer0_outputs(3707)));
    layer1_outputs(9195) <= layer0_outputs(4092);
    layer1_outputs(9196) <= (layer0_outputs(6292)) xor (layer0_outputs(301));
    layer1_outputs(9197) <= not(layer0_outputs(3943)) or (layer0_outputs(7697));
    layer1_outputs(9198) <= not(layer0_outputs(4151));
    layer1_outputs(9199) <= not(layer0_outputs(766));
    layer1_outputs(9200) <= not((layer0_outputs(80)) or (layer0_outputs(1222)));
    layer1_outputs(9201) <= layer0_outputs(2138);
    layer1_outputs(9202) <= (layer0_outputs(10084)) xor (layer0_outputs(8192));
    layer1_outputs(9203) <= not(layer0_outputs(3334));
    layer1_outputs(9204) <= layer0_outputs(276);
    layer1_outputs(9205) <= (layer0_outputs(2225)) and not (layer0_outputs(7908));
    layer1_outputs(9206) <= not(layer0_outputs(4208)) or (layer0_outputs(6205));
    layer1_outputs(9207) <= not((layer0_outputs(1728)) xor (layer0_outputs(2783)));
    layer1_outputs(9208) <= not(layer0_outputs(10109)) or (layer0_outputs(7272));
    layer1_outputs(9209) <= layer0_outputs(1410);
    layer1_outputs(9210) <= not(layer0_outputs(9328)) or (layer0_outputs(8551));
    layer1_outputs(9211) <= not((layer0_outputs(1305)) or (layer0_outputs(7420)));
    layer1_outputs(9212) <= not(layer0_outputs(3236));
    layer1_outputs(9213) <= not((layer0_outputs(3539)) xor (layer0_outputs(4936)));
    layer1_outputs(9214) <= '0';
    layer1_outputs(9215) <= not(layer0_outputs(5535));
    layer1_outputs(9216) <= not((layer0_outputs(5843)) or (layer0_outputs(2688)));
    layer1_outputs(9217) <= layer0_outputs(8513);
    layer1_outputs(9218) <= layer0_outputs(3234);
    layer1_outputs(9219) <= layer0_outputs(6006);
    layer1_outputs(9220) <= not(layer0_outputs(5594));
    layer1_outputs(9221) <= (layer0_outputs(886)) or (layer0_outputs(2239));
    layer1_outputs(9222) <= not(layer0_outputs(7154)) or (layer0_outputs(4868));
    layer1_outputs(9223) <= (layer0_outputs(2087)) and not (layer0_outputs(8120));
    layer1_outputs(9224) <= layer0_outputs(2459);
    layer1_outputs(9225) <= (layer0_outputs(9148)) and not (layer0_outputs(4768));
    layer1_outputs(9226) <= (layer0_outputs(9648)) and not (layer0_outputs(4066));
    layer1_outputs(9227) <= not((layer0_outputs(8440)) or (layer0_outputs(3868)));
    layer1_outputs(9228) <= layer0_outputs(1948);
    layer1_outputs(9229) <= (layer0_outputs(532)) xor (layer0_outputs(5221));
    layer1_outputs(9230) <= not((layer0_outputs(4200)) and (layer0_outputs(1901)));
    layer1_outputs(9231) <= not(layer0_outputs(2362)) or (layer0_outputs(4760));
    layer1_outputs(9232) <= not(layer0_outputs(8681));
    layer1_outputs(9233) <= layer0_outputs(7743);
    layer1_outputs(9234) <= not(layer0_outputs(8782));
    layer1_outputs(9235) <= layer0_outputs(9831);
    layer1_outputs(9236) <= not((layer0_outputs(2747)) or (layer0_outputs(6495)));
    layer1_outputs(9237) <= not(layer0_outputs(1712)) or (layer0_outputs(4513));
    layer1_outputs(9238) <= (layer0_outputs(8694)) and not (layer0_outputs(431));
    layer1_outputs(9239) <= not((layer0_outputs(8312)) and (layer0_outputs(6288)));
    layer1_outputs(9240) <= not(layer0_outputs(7629));
    layer1_outputs(9241) <= not(layer0_outputs(3981));
    layer1_outputs(9242) <= not(layer0_outputs(2474));
    layer1_outputs(9243) <= (layer0_outputs(4446)) xor (layer0_outputs(6435));
    layer1_outputs(9244) <= not(layer0_outputs(7241));
    layer1_outputs(9245) <= (layer0_outputs(6415)) or (layer0_outputs(4541));
    layer1_outputs(9246) <= (layer0_outputs(7750)) xor (layer0_outputs(6195));
    layer1_outputs(9247) <= (layer0_outputs(4363)) xor (layer0_outputs(156));
    layer1_outputs(9248) <= not(layer0_outputs(3032));
    layer1_outputs(9249) <= (layer0_outputs(9967)) xor (layer0_outputs(7561));
    layer1_outputs(9250) <= not(layer0_outputs(5211)) or (layer0_outputs(10192));
    layer1_outputs(9251) <= not(layer0_outputs(9004));
    layer1_outputs(9252) <= (layer0_outputs(3131)) and not (layer0_outputs(2301));
    layer1_outputs(9253) <= (layer0_outputs(7164)) and not (layer0_outputs(9564));
    layer1_outputs(9254) <= not(layer0_outputs(1288));
    layer1_outputs(9255) <= not(layer0_outputs(3338));
    layer1_outputs(9256) <= (layer0_outputs(2958)) and not (layer0_outputs(7647));
    layer1_outputs(9257) <= not(layer0_outputs(7838));
    layer1_outputs(9258) <= not(layer0_outputs(4102)) or (layer0_outputs(8228));
    layer1_outputs(9259) <= not((layer0_outputs(3720)) or (layer0_outputs(8101)));
    layer1_outputs(9260) <= layer0_outputs(7409);
    layer1_outputs(9261) <= not(layer0_outputs(4611));
    layer1_outputs(9262) <= not(layer0_outputs(3848)) or (layer0_outputs(7872));
    layer1_outputs(9263) <= (layer0_outputs(3342)) and not (layer0_outputs(5974));
    layer1_outputs(9264) <= not(layer0_outputs(6325));
    layer1_outputs(9265) <= not(layer0_outputs(5753)) or (layer0_outputs(2840));
    layer1_outputs(9266) <= layer0_outputs(9713);
    layer1_outputs(9267) <= not(layer0_outputs(8103));
    layer1_outputs(9268) <= (layer0_outputs(1537)) xor (layer0_outputs(8102));
    layer1_outputs(9269) <= '1';
    layer1_outputs(9270) <= (layer0_outputs(3929)) and (layer0_outputs(6910));
    layer1_outputs(9271) <= not(layer0_outputs(8894));
    layer1_outputs(9272) <= (layer0_outputs(3611)) or (layer0_outputs(6309));
    layer1_outputs(9273) <= layer0_outputs(5339);
    layer1_outputs(9274) <= not(layer0_outputs(1433));
    layer1_outputs(9275) <= layer0_outputs(557);
    layer1_outputs(9276) <= not((layer0_outputs(1544)) xor (layer0_outputs(2215)));
    layer1_outputs(9277) <= not((layer0_outputs(3581)) and (layer0_outputs(6759)));
    layer1_outputs(9278) <= (layer0_outputs(6921)) and (layer0_outputs(382));
    layer1_outputs(9279) <= not(layer0_outputs(2270));
    layer1_outputs(9280) <= layer0_outputs(3628);
    layer1_outputs(9281) <= not((layer0_outputs(2780)) xor (layer0_outputs(2412)));
    layer1_outputs(9282) <= not(layer0_outputs(5736));
    layer1_outputs(9283) <= not(layer0_outputs(1453));
    layer1_outputs(9284) <= not(layer0_outputs(7467)) or (layer0_outputs(487));
    layer1_outputs(9285) <= not((layer0_outputs(4616)) and (layer0_outputs(4161)));
    layer1_outputs(9286) <= layer0_outputs(4718);
    layer1_outputs(9287) <= not((layer0_outputs(7062)) or (layer0_outputs(3800)));
    layer1_outputs(9288) <= not((layer0_outputs(115)) xor (layer0_outputs(9492)));
    layer1_outputs(9289) <= not((layer0_outputs(7736)) xor (layer0_outputs(334)));
    layer1_outputs(9290) <= layer0_outputs(9094);
    layer1_outputs(9291) <= (layer0_outputs(5400)) and not (layer0_outputs(5160));
    layer1_outputs(9292) <= not((layer0_outputs(2470)) xor (layer0_outputs(8525)));
    layer1_outputs(9293) <= not(layer0_outputs(9354));
    layer1_outputs(9294) <= (layer0_outputs(6079)) and not (layer0_outputs(5267));
    layer1_outputs(9295) <= layer0_outputs(4994);
    layer1_outputs(9296) <= (layer0_outputs(2711)) or (layer0_outputs(3880));
    layer1_outputs(9297) <= (layer0_outputs(3922)) or (layer0_outputs(2980));
    layer1_outputs(9298) <= (layer0_outputs(10199)) or (layer0_outputs(2222));
    layer1_outputs(9299) <= not((layer0_outputs(2770)) xor (layer0_outputs(10213)));
    layer1_outputs(9300) <= not(layer0_outputs(5742));
    layer1_outputs(9301) <= not(layer0_outputs(3494));
    layer1_outputs(9302) <= not(layer0_outputs(7756));
    layer1_outputs(9303) <= not(layer0_outputs(4817)) or (layer0_outputs(9149));
    layer1_outputs(9304) <= not(layer0_outputs(9380));
    layer1_outputs(9305) <= layer0_outputs(6309);
    layer1_outputs(9306) <= not(layer0_outputs(9027));
    layer1_outputs(9307) <= (layer0_outputs(7907)) and not (layer0_outputs(4662));
    layer1_outputs(9308) <= not(layer0_outputs(8256)) or (layer0_outputs(7761));
    layer1_outputs(9309) <= layer0_outputs(9617);
    layer1_outputs(9310) <= not((layer0_outputs(8862)) xor (layer0_outputs(5497)));
    layer1_outputs(9311) <= not(layer0_outputs(9916));
    layer1_outputs(9312) <= (layer0_outputs(755)) or (layer0_outputs(9392));
    layer1_outputs(9313) <= not((layer0_outputs(2010)) and (layer0_outputs(55)));
    layer1_outputs(9314) <= layer0_outputs(4026);
    layer1_outputs(9315) <= (layer0_outputs(5615)) and not (layer0_outputs(3256));
    layer1_outputs(9316) <= '0';
    layer1_outputs(9317) <= (layer0_outputs(2684)) and not (layer0_outputs(7951));
    layer1_outputs(9318) <= not(layer0_outputs(384));
    layer1_outputs(9319) <= (layer0_outputs(1531)) and (layer0_outputs(10131));
    layer1_outputs(9320) <= (layer0_outputs(2668)) and not (layer0_outputs(9955));
    layer1_outputs(9321) <= (layer0_outputs(6130)) xor (layer0_outputs(5976));
    layer1_outputs(9322) <= (layer0_outputs(1001)) and (layer0_outputs(4306));
    layer1_outputs(9323) <= layer0_outputs(6905);
    layer1_outputs(9324) <= (layer0_outputs(5129)) and not (layer0_outputs(1071));
    layer1_outputs(9325) <= layer0_outputs(9225);
    layer1_outputs(9326) <= (layer0_outputs(2694)) or (layer0_outputs(3710));
    layer1_outputs(9327) <= (layer0_outputs(9920)) and (layer0_outputs(4936));
    layer1_outputs(9328) <= not(layer0_outputs(730)) or (layer0_outputs(9839));
    layer1_outputs(9329) <= (layer0_outputs(1402)) and not (layer0_outputs(2564));
    layer1_outputs(9330) <= (layer0_outputs(9895)) or (layer0_outputs(8381));
    layer1_outputs(9331) <= (layer0_outputs(4566)) or (layer0_outputs(354));
    layer1_outputs(9332) <= not(layer0_outputs(10097));
    layer1_outputs(9333) <= not((layer0_outputs(5910)) or (layer0_outputs(8366)));
    layer1_outputs(9334) <= (layer0_outputs(7399)) and not (layer0_outputs(9545));
    layer1_outputs(9335) <= layer0_outputs(4317);
    layer1_outputs(9336) <= (layer0_outputs(2704)) and not (layer0_outputs(58));
    layer1_outputs(9337) <= layer0_outputs(5487);
    layer1_outputs(9338) <= layer0_outputs(4711);
    layer1_outputs(9339) <= not((layer0_outputs(2040)) and (layer0_outputs(9990)));
    layer1_outputs(9340) <= (layer0_outputs(2518)) and not (layer0_outputs(5533));
    layer1_outputs(9341) <= not((layer0_outputs(6588)) or (layer0_outputs(7872)));
    layer1_outputs(9342) <= not(layer0_outputs(3533));
    layer1_outputs(9343) <= layer0_outputs(1246);
    layer1_outputs(9344) <= not((layer0_outputs(4297)) xor (layer0_outputs(8370)));
    layer1_outputs(9345) <= layer0_outputs(6584);
    layer1_outputs(9346) <= not(layer0_outputs(858));
    layer1_outputs(9347) <= (layer0_outputs(2782)) and not (layer0_outputs(8051));
    layer1_outputs(9348) <= (layer0_outputs(9773)) and not (layer0_outputs(5833));
    layer1_outputs(9349) <= not((layer0_outputs(1156)) and (layer0_outputs(451)));
    layer1_outputs(9350) <= layer0_outputs(5571);
    layer1_outputs(9351) <= not((layer0_outputs(759)) xor (layer0_outputs(7813)));
    layer1_outputs(9352) <= not(layer0_outputs(24));
    layer1_outputs(9353) <= layer0_outputs(4651);
    layer1_outputs(9354) <= not(layer0_outputs(4242));
    layer1_outputs(9355) <= layer0_outputs(3756);
    layer1_outputs(9356) <= not((layer0_outputs(7591)) or (layer0_outputs(1200)));
    layer1_outputs(9357) <= not((layer0_outputs(6343)) or (layer0_outputs(2976)));
    layer1_outputs(9358) <= not((layer0_outputs(3924)) or (layer0_outputs(8010)));
    layer1_outputs(9359) <= not(layer0_outputs(1473)) or (layer0_outputs(6767));
    layer1_outputs(9360) <= not((layer0_outputs(6916)) xor (layer0_outputs(3392)));
    layer1_outputs(9361) <= layer0_outputs(6231);
    layer1_outputs(9362) <= not(layer0_outputs(1915));
    layer1_outputs(9363) <= layer0_outputs(7309);
    layer1_outputs(9364) <= not(layer0_outputs(8960)) or (layer0_outputs(6204));
    layer1_outputs(9365) <= not(layer0_outputs(7721));
    layer1_outputs(9366) <= (layer0_outputs(3688)) and not (layer0_outputs(9451));
    layer1_outputs(9367) <= (layer0_outputs(9060)) or (layer0_outputs(1294));
    layer1_outputs(9368) <= not(layer0_outputs(5282));
    layer1_outputs(9369) <= not(layer0_outputs(1865)) or (layer0_outputs(6492));
    layer1_outputs(9370) <= layer0_outputs(4610);
    layer1_outputs(9371) <= not(layer0_outputs(62));
    layer1_outputs(9372) <= not(layer0_outputs(3601));
    layer1_outputs(9373) <= not(layer0_outputs(6811));
    layer1_outputs(9374) <= layer0_outputs(8767);
    layer1_outputs(9375) <= (layer0_outputs(7198)) or (layer0_outputs(169));
    layer1_outputs(9376) <= (layer0_outputs(3175)) and not (layer0_outputs(3804));
    layer1_outputs(9377) <= not(layer0_outputs(7622)) or (layer0_outputs(10137));
    layer1_outputs(9378) <= not(layer0_outputs(2884));
    layer1_outputs(9379) <= not(layer0_outputs(4617));
    layer1_outputs(9380) <= not(layer0_outputs(7625)) or (layer0_outputs(3358));
    layer1_outputs(9381) <= not(layer0_outputs(3613));
    layer1_outputs(9382) <= layer0_outputs(6518);
    layer1_outputs(9383) <= (layer0_outputs(6050)) or (layer0_outputs(3931));
    layer1_outputs(9384) <= not((layer0_outputs(4580)) xor (layer0_outputs(866)));
    layer1_outputs(9385) <= (layer0_outputs(3292)) and not (layer0_outputs(3496));
    layer1_outputs(9386) <= (layer0_outputs(1340)) and (layer0_outputs(9969));
    layer1_outputs(9387) <= layer0_outputs(6835);
    layer1_outputs(9388) <= layer0_outputs(2979);
    layer1_outputs(9389) <= (layer0_outputs(6215)) or (layer0_outputs(9926));
    layer1_outputs(9390) <= (layer0_outputs(6358)) xor (layer0_outputs(1266));
    layer1_outputs(9391) <= not(layer0_outputs(7726));
    layer1_outputs(9392) <= (layer0_outputs(520)) and (layer0_outputs(6892));
    layer1_outputs(9393) <= layer0_outputs(4019);
    layer1_outputs(9394) <= not(layer0_outputs(3293));
    layer1_outputs(9395) <= not(layer0_outputs(7973));
    layer1_outputs(9396) <= (layer0_outputs(6725)) xor (layer0_outputs(8380));
    layer1_outputs(9397) <= layer0_outputs(50);
    layer1_outputs(9398) <= not(layer0_outputs(437));
    layer1_outputs(9399) <= (layer0_outputs(3567)) and not (layer0_outputs(9800));
    layer1_outputs(9400) <= not((layer0_outputs(8053)) and (layer0_outputs(4377)));
    layer1_outputs(9401) <= not((layer0_outputs(5280)) or (layer0_outputs(247)));
    layer1_outputs(9402) <= (layer0_outputs(94)) or (layer0_outputs(8234));
    layer1_outputs(9403) <= (layer0_outputs(9608)) and not (layer0_outputs(7856));
    layer1_outputs(9404) <= not(layer0_outputs(9827));
    layer1_outputs(9405) <= not((layer0_outputs(6312)) and (layer0_outputs(4397)));
    layer1_outputs(9406) <= not(layer0_outputs(3882));
    layer1_outputs(9407) <= layer0_outputs(617);
    layer1_outputs(9408) <= not(layer0_outputs(8084));
    layer1_outputs(9409) <= layer0_outputs(8957);
    layer1_outputs(9410) <= (layer0_outputs(3459)) and not (layer0_outputs(3002));
    layer1_outputs(9411) <= not((layer0_outputs(7193)) xor (layer0_outputs(4149)));
    layer1_outputs(9412) <= not(layer0_outputs(5968));
    layer1_outputs(9413) <= (layer0_outputs(24)) or (layer0_outputs(3781));
    layer1_outputs(9414) <= layer0_outputs(1670);
    layer1_outputs(9415) <= not(layer0_outputs(3143));
    layer1_outputs(9416) <= not(layer0_outputs(4629));
    layer1_outputs(9417) <= layer0_outputs(9799);
    layer1_outputs(9418) <= not((layer0_outputs(10055)) and (layer0_outputs(6814)));
    layer1_outputs(9419) <= not(layer0_outputs(6350));
    layer1_outputs(9420) <= not((layer0_outputs(9062)) and (layer0_outputs(7227)));
    layer1_outputs(9421) <= not(layer0_outputs(6369)) or (layer0_outputs(1947));
    layer1_outputs(9422) <= layer0_outputs(7893);
    layer1_outputs(9423) <= not((layer0_outputs(7678)) and (layer0_outputs(1321)));
    layer1_outputs(9424) <= (layer0_outputs(2623)) and not (layer0_outputs(364));
    layer1_outputs(9425) <= not((layer0_outputs(8068)) or (layer0_outputs(6374)));
    layer1_outputs(9426) <= not(layer0_outputs(7796));
    layer1_outputs(9427) <= not(layer0_outputs(2064));
    layer1_outputs(9428) <= '0';
    layer1_outputs(9429) <= layer0_outputs(8303);
    layer1_outputs(9430) <= (layer0_outputs(6141)) and not (layer0_outputs(9092));
    layer1_outputs(9431) <= not((layer0_outputs(3171)) and (layer0_outputs(8235)));
    layer1_outputs(9432) <= not((layer0_outputs(3213)) and (layer0_outputs(6889)));
    layer1_outputs(9433) <= not(layer0_outputs(2757));
    layer1_outputs(9434) <= not((layer0_outputs(9134)) or (layer0_outputs(8699)));
    layer1_outputs(9435) <= (layer0_outputs(4891)) or (layer0_outputs(7993));
    layer1_outputs(9436) <= layer0_outputs(7530);
    layer1_outputs(9437) <= (layer0_outputs(6245)) and not (layer0_outputs(2951));
    layer1_outputs(9438) <= not(layer0_outputs(7249));
    layer1_outputs(9439) <= not((layer0_outputs(3241)) and (layer0_outputs(4817)));
    layer1_outputs(9440) <= not(layer0_outputs(5529));
    layer1_outputs(9441) <= (layer0_outputs(3637)) and not (layer0_outputs(3369));
    layer1_outputs(9442) <= (layer0_outputs(5577)) xor (layer0_outputs(7768));
    layer1_outputs(9443) <= not((layer0_outputs(8954)) and (layer0_outputs(10048)));
    layer1_outputs(9444) <= (layer0_outputs(6716)) and (layer0_outputs(7087));
    layer1_outputs(9445) <= not((layer0_outputs(4973)) or (layer0_outputs(3284)));
    layer1_outputs(9446) <= '0';
    layer1_outputs(9447) <= not(layer0_outputs(5114));
    layer1_outputs(9448) <= layer0_outputs(142);
    layer1_outputs(9449) <= not(layer0_outputs(1561));
    layer1_outputs(9450) <= not(layer0_outputs(9064));
    layer1_outputs(9451) <= not((layer0_outputs(884)) xor (layer0_outputs(4297)));
    layer1_outputs(9452) <= not(layer0_outputs(8190)) or (layer0_outputs(949));
    layer1_outputs(9453) <= not(layer0_outputs(2421));
    layer1_outputs(9454) <= layer0_outputs(8225);
    layer1_outputs(9455) <= not(layer0_outputs(9968));
    layer1_outputs(9456) <= not((layer0_outputs(6511)) xor (layer0_outputs(9563)));
    layer1_outputs(9457) <= not(layer0_outputs(525));
    layer1_outputs(9458) <= (layer0_outputs(9102)) and not (layer0_outputs(7982));
    layer1_outputs(9459) <= not((layer0_outputs(4003)) xor (layer0_outputs(6217)));
    layer1_outputs(9460) <= (layer0_outputs(7040)) or (layer0_outputs(8421));
    layer1_outputs(9461) <= (layer0_outputs(646)) and not (layer0_outputs(540));
    layer1_outputs(9462) <= not(layer0_outputs(3378)) or (layer0_outputs(6172));
    layer1_outputs(9463) <= not(layer0_outputs(6620)) or (layer0_outputs(8724));
    layer1_outputs(9464) <= layer0_outputs(4289);
    layer1_outputs(9465) <= not((layer0_outputs(3588)) or (layer0_outputs(733)));
    layer1_outputs(9466) <= not(layer0_outputs(4548));
    layer1_outputs(9467) <= not((layer0_outputs(9977)) or (layer0_outputs(8613)));
    layer1_outputs(9468) <= (layer0_outputs(7715)) or (layer0_outputs(3337));
    layer1_outputs(9469) <= (layer0_outputs(8205)) and not (layer0_outputs(5627));
    layer1_outputs(9470) <= not((layer0_outputs(5994)) xor (layer0_outputs(208)));
    layer1_outputs(9471) <= not(layer0_outputs(8444));
    layer1_outputs(9472) <= (layer0_outputs(1898)) and not (layer0_outputs(3212));
    layer1_outputs(9473) <= not(layer0_outputs(6728));
    layer1_outputs(9474) <= layer0_outputs(1536);
    layer1_outputs(9475) <= not((layer0_outputs(2589)) and (layer0_outputs(8303)));
    layer1_outputs(9476) <= not(layer0_outputs(8229));
    layer1_outputs(9477) <= layer0_outputs(1515);
    layer1_outputs(9478) <= (layer0_outputs(4509)) or (layer0_outputs(9930));
    layer1_outputs(9479) <= (layer0_outputs(6054)) and not (layer0_outputs(9954));
    layer1_outputs(9480) <= not((layer0_outputs(5517)) or (layer0_outputs(10014)));
    layer1_outputs(9481) <= not(layer0_outputs(7821));
    layer1_outputs(9482) <= (layer0_outputs(5578)) xor (layer0_outputs(2745));
    layer1_outputs(9483) <= (layer0_outputs(6599)) and (layer0_outputs(3465));
    layer1_outputs(9484) <= not((layer0_outputs(1542)) or (layer0_outputs(8288)));
    layer1_outputs(9485) <= (layer0_outputs(5212)) and not (layer0_outputs(324));
    layer1_outputs(9486) <= layer0_outputs(3735);
    layer1_outputs(9487) <= (layer0_outputs(3906)) or (layer0_outputs(9308));
    layer1_outputs(9488) <= not(layer0_outputs(4995));
    layer1_outputs(9489) <= (layer0_outputs(3690)) and not (layer0_outputs(2453));
    layer1_outputs(9490) <= (layer0_outputs(5098)) and not (layer0_outputs(9695));
    layer1_outputs(9491) <= (layer0_outputs(3759)) and not (layer0_outputs(5819));
    layer1_outputs(9492) <= layer0_outputs(5791);
    layer1_outputs(9493) <= not(layer0_outputs(7875));
    layer1_outputs(9494) <= not(layer0_outputs(6253)) or (layer0_outputs(9208));
    layer1_outputs(9495) <= (layer0_outputs(64)) and not (layer0_outputs(1033));
    layer1_outputs(9496) <= (layer0_outputs(8926)) and not (layer0_outputs(1500));
    layer1_outputs(9497) <= (layer0_outputs(2596)) and not (layer0_outputs(7338));
    layer1_outputs(9498) <= not((layer0_outputs(6335)) and (layer0_outputs(1272)));
    layer1_outputs(9499) <= not(layer0_outputs(5003));
    layer1_outputs(9500) <= layer0_outputs(4074);
    layer1_outputs(9501) <= (layer0_outputs(635)) and not (layer0_outputs(4114));
    layer1_outputs(9502) <= (layer0_outputs(6568)) and (layer0_outputs(960));
    layer1_outputs(9503) <= not(layer0_outputs(6551));
    layer1_outputs(9504) <= (layer0_outputs(9509)) and not (layer0_outputs(6218));
    layer1_outputs(9505) <= not(layer0_outputs(4001)) or (layer0_outputs(2751));
    layer1_outputs(9506) <= not(layer0_outputs(3158));
    layer1_outputs(9507) <= layer0_outputs(493);
    layer1_outputs(9508) <= not((layer0_outputs(7871)) or (layer0_outputs(7941)));
    layer1_outputs(9509) <= layer0_outputs(5647);
    layer1_outputs(9510) <= layer0_outputs(6597);
    layer1_outputs(9511) <= layer0_outputs(6969);
    layer1_outputs(9512) <= (layer0_outputs(4367)) and (layer0_outputs(3689));
    layer1_outputs(9513) <= layer0_outputs(9180);
    layer1_outputs(9514) <= '0';
    layer1_outputs(9515) <= layer0_outputs(9791);
    layer1_outputs(9516) <= not((layer0_outputs(5845)) xor (layer0_outputs(7352)));
    layer1_outputs(9517) <= (layer0_outputs(1770)) and not (layer0_outputs(617));
    layer1_outputs(9518) <= (layer0_outputs(2004)) and (layer0_outputs(9251));
    layer1_outputs(9519) <= (layer0_outputs(8087)) and not (layer0_outputs(9055));
    layer1_outputs(9520) <= not((layer0_outputs(713)) xor (layer0_outputs(8988)));
    layer1_outputs(9521) <= not(layer0_outputs(4848));
    layer1_outputs(9522) <= layer0_outputs(9275);
    layer1_outputs(9523) <= layer0_outputs(9422);
    layer1_outputs(9524) <= not(layer0_outputs(5615));
    layer1_outputs(9525) <= not(layer0_outputs(22));
    layer1_outputs(9526) <= layer0_outputs(2343);
    layer1_outputs(9527) <= not(layer0_outputs(6331));
    layer1_outputs(9528) <= (layer0_outputs(9716)) and not (layer0_outputs(1007));
    layer1_outputs(9529) <= not(layer0_outputs(5898)) or (layer0_outputs(6624));
    layer1_outputs(9530) <= layer0_outputs(5936);
    layer1_outputs(9531) <= not(layer0_outputs(352));
    layer1_outputs(9532) <= not(layer0_outputs(10202)) or (layer0_outputs(3061));
    layer1_outputs(9533) <= not(layer0_outputs(3788)) or (layer0_outputs(6866));
    layer1_outputs(9534) <= not(layer0_outputs(6755)) or (layer0_outputs(9224));
    layer1_outputs(9535) <= (layer0_outputs(9141)) xor (layer0_outputs(8689));
    layer1_outputs(9536) <= not((layer0_outputs(4798)) xor (layer0_outputs(8301)));
    layer1_outputs(9537) <= layer0_outputs(9572);
    layer1_outputs(9538) <= '0';
    layer1_outputs(9539) <= (layer0_outputs(10098)) and not (layer0_outputs(2275));
    layer1_outputs(9540) <= layer0_outputs(4709);
    layer1_outputs(9541) <= (layer0_outputs(3767)) and not (layer0_outputs(1450));
    layer1_outputs(9542) <= not((layer0_outputs(6077)) and (layer0_outputs(9055)));
    layer1_outputs(9543) <= not((layer0_outputs(1224)) and (layer0_outputs(6956)));
    layer1_outputs(9544) <= layer0_outputs(7307);
    layer1_outputs(9545) <= not(layer0_outputs(5548)) or (layer0_outputs(3642));
    layer1_outputs(9546) <= not((layer0_outputs(6837)) and (layer0_outputs(7034)));
    layer1_outputs(9547) <= not(layer0_outputs(8786));
    layer1_outputs(9548) <= not((layer0_outputs(1199)) and (layer0_outputs(7335)));
    layer1_outputs(9549) <= (layer0_outputs(7502)) and not (layer0_outputs(7649));
    layer1_outputs(9550) <= not((layer0_outputs(6615)) or (layer0_outputs(1125)));
    layer1_outputs(9551) <= layer0_outputs(4319);
    layer1_outputs(9552) <= not(layer0_outputs(9726));
    layer1_outputs(9553) <= not((layer0_outputs(4184)) or (layer0_outputs(3801)));
    layer1_outputs(9554) <= layer0_outputs(4596);
    layer1_outputs(9555) <= '0';
    layer1_outputs(9556) <= not((layer0_outputs(8959)) xor (layer0_outputs(4142)));
    layer1_outputs(9557) <= layer0_outputs(2641);
    layer1_outputs(9558) <= not(layer0_outputs(1788));
    layer1_outputs(9559) <= (layer0_outputs(10036)) and not (layer0_outputs(7531));
    layer1_outputs(9560) <= (layer0_outputs(7524)) and (layer0_outputs(3774));
    layer1_outputs(9561) <= not(layer0_outputs(7116));
    layer1_outputs(9562) <= (layer0_outputs(6140)) and (layer0_outputs(727));
    layer1_outputs(9563) <= layer0_outputs(7140);
    layer1_outputs(9564) <= layer0_outputs(9232);
    layer1_outputs(9565) <= (layer0_outputs(8150)) and (layer0_outputs(9829));
    layer1_outputs(9566) <= not((layer0_outputs(8716)) and (layer0_outputs(269)));
    layer1_outputs(9567) <= (layer0_outputs(8895)) or (layer0_outputs(2437));
    layer1_outputs(9568) <= (layer0_outputs(8556)) or (layer0_outputs(9357));
    layer1_outputs(9569) <= (layer0_outputs(2693)) and not (layer0_outputs(2702));
    layer1_outputs(9570) <= (layer0_outputs(5566)) or (layer0_outputs(8570));
    layer1_outputs(9571) <= layer0_outputs(6085);
    layer1_outputs(9572) <= not(layer0_outputs(4346)) or (layer0_outputs(6493));
    layer1_outputs(9573) <= not((layer0_outputs(9074)) or (layer0_outputs(9292)));
    layer1_outputs(9574) <= (layer0_outputs(8245)) or (layer0_outputs(8336));
    layer1_outputs(9575) <= (layer0_outputs(1333)) and (layer0_outputs(1950));
    layer1_outputs(9576) <= layer0_outputs(2195);
    layer1_outputs(9577) <= layer0_outputs(9851);
    layer1_outputs(9578) <= not((layer0_outputs(2407)) and (layer0_outputs(8131)));
    layer1_outputs(9579) <= not(layer0_outputs(7016));
    layer1_outputs(9580) <= not(layer0_outputs(5760));
    layer1_outputs(9581) <= (layer0_outputs(2744)) or (layer0_outputs(4099));
    layer1_outputs(9582) <= not(layer0_outputs(5056));
    layer1_outputs(9583) <= (layer0_outputs(4752)) and (layer0_outputs(1503));
    layer1_outputs(9584) <= not(layer0_outputs(1238));
    layer1_outputs(9585) <= (layer0_outputs(8760)) or (layer0_outputs(5300));
    layer1_outputs(9586) <= not(layer0_outputs(2089));
    layer1_outputs(9587) <= layer0_outputs(4254);
    layer1_outputs(9588) <= (layer0_outputs(3785)) and not (layer0_outputs(6967));
    layer1_outputs(9589) <= not(layer0_outputs(6816)) or (layer0_outputs(4240));
    layer1_outputs(9590) <= layer0_outputs(9932);
    layer1_outputs(9591) <= (layer0_outputs(4147)) or (layer0_outputs(5246));
    layer1_outputs(9592) <= layer0_outputs(9594);
    layer1_outputs(9593) <= not(layer0_outputs(4650));
    layer1_outputs(9594) <= not(layer0_outputs(3026));
    layer1_outputs(9595) <= not(layer0_outputs(3593)) or (layer0_outputs(3875));
    layer1_outputs(9596) <= layer0_outputs(1207);
    layer1_outputs(9597) <= not(layer0_outputs(1403)) or (layer0_outputs(2136));
    layer1_outputs(9598) <= layer0_outputs(7020);
    layer1_outputs(9599) <= not(layer0_outputs(8565)) or (layer0_outputs(4557));
    layer1_outputs(9600) <= layer0_outputs(4481);
    layer1_outputs(9601) <= not(layer0_outputs(5514)) or (layer0_outputs(3708));
    layer1_outputs(9602) <= layer0_outputs(3207);
    layer1_outputs(9603) <= (layer0_outputs(5022)) xor (layer0_outputs(537));
    layer1_outputs(9604) <= not(layer0_outputs(6110)) or (layer0_outputs(9961));
    layer1_outputs(9605) <= (layer0_outputs(1284)) and not (layer0_outputs(4247));
    layer1_outputs(9606) <= not((layer0_outputs(3138)) or (layer0_outputs(2750)));
    layer1_outputs(9607) <= not((layer0_outputs(3042)) xor (layer0_outputs(3534)));
    layer1_outputs(9608) <= not((layer0_outputs(6486)) and (layer0_outputs(1531)));
    layer1_outputs(9609) <= not((layer0_outputs(8913)) or (layer0_outputs(3594)));
    layer1_outputs(9610) <= not(layer0_outputs(2585));
    layer1_outputs(9611) <= (layer0_outputs(9243)) or (layer0_outputs(89));
    layer1_outputs(9612) <= not(layer0_outputs(2370)) or (layer0_outputs(8619));
    layer1_outputs(9613) <= (layer0_outputs(3055)) and not (layer0_outputs(8));
    layer1_outputs(9614) <= (layer0_outputs(6032)) xor (layer0_outputs(1387));
    layer1_outputs(9615) <= layer0_outputs(3383);
    layer1_outputs(9616) <= layer0_outputs(6151);
    layer1_outputs(9617) <= (layer0_outputs(4922)) and not (layer0_outputs(2920));
    layer1_outputs(9618) <= not((layer0_outputs(9569)) and (layer0_outputs(4071)));
    layer1_outputs(9619) <= layer0_outputs(4528);
    layer1_outputs(9620) <= not((layer0_outputs(1198)) xor (layer0_outputs(5718)));
    layer1_outputs(9621) <= layer0_outputs(201);
    layer1_outputs(9622) <= not(layer0_outputs(1956)) or (layer0_outputs(2317));
    layer1_outputs(9623) <= not(layer0_outputs(2912));
    layer1_outputs(9624) <= not(layer0_outputs(4457)) or (layer0_outputs(1565));
    layer1_outputs(9625) <= layer0_outputs(170);
    layer1_outputs(9626) <= (layer0_outputs(5959)) and not (layer0_outputs(7208));
    layer1_outputs(9627) <= (layer0_outputs(3697)) and not (layer0_outputs(735));
    layer1_outputs(9628) <= (layer0_outputs(8844)) and (layer0_outputs(3624));
    layer1_outputs(9629) <= (layer0_outputs(2831)) and not (layer0_outputs(2914));
    layer1_outputs(9630) <= layer0_outputs(6307);
    layer1_outputs(9631) <= (layer0_outputs(45)) or (layer0_outputs(3079));
    layer1_outputs(9632) <= layer0_outputs(8591);
    layer1_outputs(9633) <= '0';
    layer1_outputs(9634) <= (layer0_outputs(8743)) and not (layer0_outputs(8195));
    layer1_outputs(9635) <= layer0_outputs(5334);
    layer1_outputs(9636) <= not(layer0_outputs(9091)) or (layer0_outputs(9303));
    layer1_outputs(9637) <= not((layer0_outputs(5466)) and (layer0_outputs(8995)));
    layer1_outputs(9638) <= (layer0_outputs(1308)) xor (layer0_outputs(4846));
    layer1_outputs(9639) <= (layer0_outputs(3946)) and (layer0_outputs(4107));
    layer1_outputs(9640) <= not(layer0_outputs(4313)) or (layer0_outputs(6634));
    layer1_outputs(9641) <= layer0_outputs(571);
    layer1_outputs(9642) <= not((layer0_outputs(4147)) or (layer0_outputs(190)));
    layer1_outputs(9643) <= layer0_outputs(5732);
    layer1_outputs(9644) <= not(layer0_outputs(8857)) or (layer0_outputs(9376));
    layer1_outputs(9645) <= not((layer0_outputs(3699)) and (layer0_outputs(4866)));
    layer1_outputs(9646) <= not((layer0_outputs(4173)) and (layer0_outputs(7339)));
    layer1_outputs(9647) <= layer0_outputs(4036);
    layer1_outputs(9648) <= not((layer0_outputs(7212)) xor (layer0_outputs(4889)));
    layer1_outputs(9649) <= (layer0_outputs(671)) or (layer0_outputs(6632));
    layer1_outputs(9650) <= not(layer0_outputs(9891));
    layer1_outputs(9651) <= not(layer0_outputs(5322));
    layer1_outputs(9652) <= not(layer0_outputs(7857)) or (layer0_outputs(3830));
    layer1_outputs(9653) <= not(layer0_outputs(6898));
    layer1_outputs(9654) <= layer0_outputs(5931);
    layer1_outputs(9655) <= layer0_outputs(9940);
    layer1_outputs(9656) <= not(layer0_outputs(8111)) or (layer0_outputs(347));
    layer1_outputs(9657) <= layer0_outputs(8382);
    layer1_outputs(9658) <= not(layer0_outputs(88));
    layer1_outputs(9659) <= (layer0_outputs(8187)) and not (layer0_outputs(6200));
    layer1_outputs(9660) <= not(layer0_outputs(5934)) or (layer0_outputs(5376));
    layer1_outputs(9661) <= (layer0_outputs(7225)) xor (layer0_outputs(2420));
    layer1_outputs(9662) <= not(layer0_outputs(3641)) or (layer0_outputs(1170));
    layer1_outputs(9663) <= (layer0_outputs(996)) and not (layer0_outputs(696));
    layer1_outputs(9664) <= not(layer0_outputs(880)) or (layer0_outputs(2134));
    layer1_outputs(9665) <= (layer0_outputs(8488)) and (layer0_outputs(8435));
    layer1_outputs(9666) <= not((layer0_outputs(5451)) or (layer0_outputs(1113)));
    layer1_outputs(9667) <= (layer0_outputs(35)) xor (layer0_outputs(8829));
    layer1_outputs(9668) <= '0';
    layer1_outputs(9669) <= (layer0_outputs(8740)) xor (layer0_outputs(10034));
    layer1_outputs(9670) <= (layer0_outputs(6158)) and (layer0_outputs(3299));
    layer1_outputs(9671) <= not(layer0_outputs(2844)) or (layer0_outputs(5595));
    layer1_outputs(9672) <= not(layer0_outputs(6963)) or (layer0_outputs(8519));
    layer1_outputs(9673) <= layer0_outputs(8825);
    layer1_outputs(9674) <= (layer0_outputs(6638)) and not (layer0_outputs(4397));
    layer1_outputs(9675) <= not((layer0_outputs(2932)) and (layer0_outputs(8322)));
    layer1_outputs(9676) <= (layer0_outputs(7033)) xor (layer0_outputs(2484));
    layer1_outputs(9677) <= (layer0_outputs(9873)) and not (layer0_outputs(4046));
    layer1_outputs(9678) <= not((layer0_outputs(2541)) or (layer0_outputs(180)));
    layer1_outputs(9679) <= not(layer0_outputs(729));
    layer1_outputs(9680) <= layer0_outputs(2380);
    layer1_outputs(9681) <= layer0_outputs(6843);
    layer1_outputs(9682) <= layer0_outputs(565);
    layer1_outputs(9683) <= '0';
    layer1_outputs(9684) <= '1';
    layer1_outputs(9685) <= not(layer0_outputs(9732));
    layer1_outputs(9686) <= (layer0_outputs(359)) and not (layer0_outputs(9336));
    layer1_outputs(9687) <= '0';
    layer1_outputs(9688) <= not(layer0_outputs(1737));
    layer1_outputs(9689) <= (layer0_outputs(7847)) and not (layer0_outputs(9027));
    layer1_outputs(9690) <= not(layer0_outputs(4211)) or (layer0_outputs(7983));
    layer1_outputs(9691) <= (layer0_outputs(3260)) xor (layer0_outputs(3635));
    layer1_outputs(9692) <= not(layer0_outputs(7412)) or (layer0_outputs(4348));
    layer1_outputs(9693) <= not(layer0_outputs(6427));
    layer1_outputs(9694) <= not(layer0_outputs(2811));
    layer1_outputs(9695) <= not(layer0_outputs(9261));
    layer1_outputs(9696) <= not(layer0_outputs(1564));
    layer1_outputs(9697) <= (layer0_outputs(7888)) xor (layer0_outputs(7188));
    layer1_outputs(9698) <= not(layer0_outputs(9070)) or (layer0_outputs(6797));
    layer1_outputs(9699) <= (layer0_outputs(3086)) or (layer0_outputs(1631));
    layer1_outputs(9700) <= layer0_outputs(8078);
    layer1_outputs(9701) <= layer0_outputs(429);
    layer1_outputs(9702) <= (layer0_outputs(1231)) and (layer0_outputs(3005));
    layer1_outputs(9703) <= (layer0_outputs(5806)) and (layer0_outputs(293));
    layer1_outputs(9704) <= (layer0_outputs(7729)) or (layer0_outputs(2497));
    layer1_outputs(9705) <= (layer0_outputs(4814)) and not (layer0_outputs(2845));
    layer1_outputs(9706) <= not((layer0_outputs(8786)) xor (layer0_outputs(7555)));
    layer1_outputs(9707) <= layer0_outputs(29);
    layer1_outputs(9708) <= (layer0_outputs(8482)) and not (layer0_outputs(5149));
    layer1_outputs(9709) <= '1';
    layer1_outputs(9710) <= layer0_outputs(5712);
    layer1_outputs(9711) <= layer0_outputs(3039);
    layer1_outputs(9712) <= (layer0_outputs(4567)) and not (layer0_outputs(1265));
    layer1_outputs(9713) <= not(layer0_outputs(1760));
    layer1_outputs(9714) <= (layer0_outputs(6000)) and (layer0_outputs(4595));
    layer1_outputs(9715) <= not((layer0_outputs(8799)) xor (layer0_outputs(1637)));
    layer1_outputs(9716) <= not(layer0_outputs(4536));
    layer1_outputs(9717) <= not(layer0_outputs(4895));
    layer1_outputs(9718) <= not(layer0_outputs(2421));
    layer1_outputs(9719) <= (layer0_outputs(3581)) xor (layer0_outputs(1517));
    layer1_outputs(9720) <= (layer0_outputs(2555)) xor (layer0_outputs(7360));
    layer1_outputs(9721) <= '1';
    layer1_outputs(9722) <= (layer0_outputs(2726)) and not (layer0_outputs(7260));
    layer1_outputs(9723) <= layer0_outputs(4424);
    layer1_outputs(9724) <= not(layer0_outputs(7069)) or (layer0_outputs(236));
    layer1_outputs(9725) <= not(layer0_outputs(5661)) or (layer0_outputs(2358));
    layer1_outputs(9726) <= not(layer0_outputs(3668));
    layer1_outputs(9727) <= (layer0_outputs(6626)) and not (layer0_outputs(1267));
    layer1_outputs(9728) <= (layer0_outputs(9826)) and (layer0_outputs(5175));
    layer1_outputs(9729) <= not(layer0_outputs(7816));
    layer1_outputs(9730) <= not((layer0_outputs(1062)) or (layer0_outputs(7689)));
    layer1_outputs(9731) <= not((layer0_outputs(933)) xor (layer0_outputs(6008)));
    layer1_outputs(9732) <= layer0_outputs(4711);
    layer1_outputs(9733) <= layer0_outputs(606);
    layer1_outputs(9734) <= not(layer0_outputs(9210)) or (layer0_outputs(747));
    layer1_outputs(9735) <= layer0_outputs(9761);
    layer1_outputs(9736) <= (layer0_outputs(5604)) and (layer0_outputs(1381));
    layer1_outputs(9737) <= not(layer0_outputs(1608));
    layer1_outputs(9738) <= not(layer0_outputs(1336));
    layer1_outputs(9739) <= '0';
    layer1_outputs(9740) <= (layer0_outputs(9543)) or (layer0_outputs(5019));
    layer1_outputs(9741) <= (layer0_outputs(216)) and (layer0_outputs(4547));
    layer1_outputs(9742) <= not(layer0_outputs(6536)) or (layer0_outputs(8757));
    layer1_outputs(9743) <= (layer0_outputs(10154)) and not (layer0_outputs(8788));
    layer1_outputs(9744) <= not((layer0_outputs(10193)) and (layer0_outputs(3422)));
    layer1_outputs(9745) <= (layer0_outputs(5919)) xor (layer0_outputs(6769));
    layer1_outputs(9746) <= (layer0_outputs(2940)) or (layer0_outputs(5320));
    layer1_outputs(9747) <= not(layer0_outputs(1412)) or (layer0_outputs(4969));
    layer1_outputs(9748) <= layer0_outputs(4660);
    layer1_outputs(9749) <= not((layer0_outputs(9201)) or (layer0_outputs(2567)));
    layer1_outputs(9750) <= not((layer0_outputs(3365)) or (layer0_outputs(8785)));
    layer1_outputs(9751) <= not(layer0_outputs(3376)) or (layer0_outputs(3394));
    layer1_outputs(9752) <= not((layer0_outputs(5137)) and (layer0_outputs(2963)));
    layer1_outputs(9753) <= layer0_outputs(8980);
    layer1_outputs(9754) <= layer0_outputs(5353);
    layer1_outputs(9755) <= not(layer0_outputs(1727));
    layer1_outputs(9756) <= (layer0_outputs(1573)) xor (layer0_outputs(4714));
    layer1_outputs(9757) <= not(layer0_outputs(3701));
    layer1_outputs(9758) <= (layer0_outputs(7332)) and not (layer0_outputs(7552));
    layer1_outputs(9759) <= not(layer0_outputs(4160));
    layer1_outputs(9760) <= layer0_outputs(10110);
    layer1_outputs(9761) <= not(layer0_outputs(7810));
    layer1_outputs(9762) <= '0';
    layer1_outputs(9763) <= layer0_outputs(7842);
    layer1_outputs(9764) <= layer0_outputs(2409);
    layer1_outputs(9765) <= layer0_outputs(3980);
    layer1_outputs(9766) <= not((layer0_outputs(223)) or (layer0_outputs(2365)));
    layer1_outputs(9767) <= not((layer0_outputs(6052)) xor (layer0_outputs(8998)));
    layer1_outputs(9768) <= (layer0_outputs(2913)) xor (layer0_outputs(8940));
    layer1_outputs(9769) <= not((layer0_outputs(7755)) xor (layer0_outputs(8121)));
    layer1_outputs(9770) <= layer0_outputs(5324);
    layer1_outputs(9771) <= not((layer0_outputs(9486)) xor (layer0_outputs(9331)));
    layer1_outputs(9772) <= not(layer0_outputs(4883)) or (layer0_outputs(4095));
    layer1_outputs(9773) <= layer0_outputs(217);
    layer1_outputs(9774) <= not(layer0_outputs(6708));
    layer1_outputs(9775) <= (layer0_outputs(2351)) and not (layer0_outputs(4545));
    layer1_outputs(9776) <= not((layer0_outputs(3789)) or (layer0_outputs(7053)));
    layer1_outputs(9777) <= (layer0_outputs(5927)) and (layer0_outputs(5244));
    layer1_outputs(9778) <= not(layer0_outputs(5465));
    layer1_outputs(9779) <= not((layer0_outputs(6416)) and (layer0_outputs(5777)));
    layer1_outputs(9780) <= layer0_outputs(9514);
    layer1_outputs(9781) <= not((layer0_outputs(7991)) or (layer0_outputs(7175)));
    layer1_outputs(9782) <= '1';
    layer1_outputs(9783) <= not((layer0_outputs(4667)) and (layer0_outputs(5902)));
    layer1_outputs(9784) <= not(layer0_outputs(1502)) or (layer0_outputs(5016));
    layer1_outputs(9785) <= '0';
    layer1_outputs(9786) <= not(layer0_outputs(1011));
    layer1_outputs(9787) <= not(layer0_outputs(3315));
    layer1_outputs(9788) <= not(layer0_outputs(2945)) or (layer0_outputs(997));
    layer1_outputs(9789) <= not(layer0_outputs(7822));
    layer1_outputs(9790) <= (layer0_outputs(7350)) and (layer0_outputs(9603));
    layer1_outputs(9791) <= not(layer0_outputs(564)) or (layer0_outputs(835));
    layer1_outputs(9792) <= (layer0_outputs(3362)) and (layer0_outputs(8550));
    layer1_outputs(9793) <= (layer0_outputs(9766)) or (layer0_outputs(7454));
    layer1_outputs(9794) <= layer0_outputs(9862);
    layer1_outputs(9795) <= not(layer0_outputs(7581));
    layer1_outputs(9796) <= not((layer0_outputs(84)) and (layer0_outputs(6245)));
    layer1_outputs(9797) <= not(layer0_outputs(5192));
    layer1_outputs(9798) <= (layer0_outputs(3952)) and not (layer0_outputs(4448));
    layer1_outputs(9799) <= not(layer0_outputs(6956));
    layer1_outputs(9800) <= (layer0_outputs(2706)) xor (layer0_outputs(6738));
    layer1_outputs(9801) <= not(layer0_outputs(4867)) or (layer0_outputs(851));
    layer1_outputs(9802) <= layer0_outputs(7395);
    layer1_outputs(9803) <= not(layer0_outputs(5876)) or (layer0_outputs(2371));
    layer1_outputs(9804) <= (layer0_outputs(2543)) and not (layer0_outputs(1693));
    layer1_outputs(9805) <= not((layer0_outputs(5294)) or (layer0_outputs(5308)));
    layer1_outputs(9806) <= not((layer0_outputs(6616)) and (layer0_outputs(1963)));
    layer1_outputs(9807) <= not((layer0_outputs(5664)) and (layer0_outputs(9862)));
    layer1_outputs(9808) <= not(layer0_outputs(2124)) or (layer0_outputs(2567));
    layer1_outputs(9809) <= '0';
    layer1_outputs(9810) <= not((layer0_outputs(3190)) xor (layer0_outputs(9775)));
    layer1_outputs(9811) <= not(layer0_outputs(1927));
    layer1_outputs(9812) <= (layer0_outputs(3060)) and not (layer0_outputs(5188));
    layer1_outputs(9813) <= not((layer0_outputs(4798)) or (layer0_outputs(9792)));
    layer1_outputs(9814) <= not((layer0_outputs(3119)) and (layer0_outputs(6859)));
    layer1_outputs(9815) <= layer0_outputs(6825);
    layer1_outputs(9816) <= not(layer0_outputs(788));
    layer1_outputs(9817) <= not(layer0_outputs(6523));
    layer1_outputs(9818) <= (layer0_outputs(3460)) and not (layer0_outputs(6801));
    layer1_outputs(9819) <= layer0_outputs(8818);
    layer1_outputs(9820) <= (layer0_outputs(9175)) or (layer0_outputs(4486));
    layer1_outputs(9821) <= not(layer0_outputs(7217));
    layer1_outputs(9822) <= (layer0_outputs(2347)) and not (layer0_outputs(3307));
    layer1_outputs(9823) <= not(layer0_outputs(3406));
    layer1_outputs(9824) <= not(layer0_outputs(5924)) or (layer0_outputs(3281));
    layer1_outputs(9825) <= (layer0_outputs(4675)) and (layer0_outputs(8839));
    layer1_outputs(9826) <= (layer0_outputs(5227)) xor (layer0_outputs(3357));
    layer1_outputs(9827) <= not((layer0_outputs(9403)) or (layer0_outputs(9616)));
    layer1_outputs(9828) <= (layer0_outputs(8796)) and not (layer0_outputs(1655));
    layer1_outputs(9829) <= not((layer0_outputs(4263)) or (layer0_outputs(5752)));
    layer1_outputs(9830) <= not(layer0_outputs(9324)) or (layer0_outputs(9309));
    layer1_outputs(9831) <= not((layer0_outputs(7488)) xor (layer0_outputs(1240)));
    layer1_outputs(9832) <= (layer0_outputs(6058)) and not (layer0_outputs(7135));
    layer1_outputs(9833) <= layer0_outputs(9937);
    layer1_outputs(9834) <= not(layer0_outputs(2267)) or (layer0_outputs(994));
    layer1_outputs(9835) <= not(layer0_outputs(3451));
    layer1_outputs(9836) <= layer0_outputs(7372);
    layer1_outputs(9837) <= not(layer0_outputs(2399)) or (layer0_outputs(1419));
    layer1_outputs(9838) <= not(layer0_outputs(556));
    layer1_outputs(9839) <= layer0_outputs(4816);
    layer1_outputs(9840) <= not((layer0_outputs(773)) and (layer0_outputs(10230)));
    layer1_outputs(9841) <= not(layer0_outputs(5709)) or (layer0_outputs(9455));
    layer1_outputs(9842) <= layer0_outputs(7746);
    layer1_outputs(9843) <= layer0_outputs(2141);
    layer1_outputs(9844) <= not(layer0_outputs(6719));
    layer1_outputs(9845) <= not(layer0_outputs(1122)) or (layer0_outputs(9724));
    layer1_outputs(9846) <= not((layer0_outputs(1529)) and (layer0_outputs(3597)));
    layer1_outputs(9847) <= not(layer0_outputs(3961));
    layer1_outputs(9848) <= not(layer0_outputs(7304)) or (layer0_outputs(1312));
    layer1_outputs(9849) <= layer0_outputs(4029);
    layer1_outputs(9850) <= not(layer0_outputs(1396));
    layer1_outputs(9851) <= not((layer0_outputs(1218)) or (layer0_outputs(2830)));
    layer1_outputs(9852) <= layer0_outputs(5719);
    layer1_outputs(9853) <= (layer0_outputs(10232)) or (layer0_outputs(746));
    layer1_outputs(9854) <= not(layer0_outputs(2982));
    layer1_outputs(9855) <= layer0_outputs(2597);
    layer1_outputs(9856) <= (layer0_outputs(2710)) xor (layer0_outputs(3526));
    layer1_outputs(9857) <= layer0_outputs(2942);
    layer1_outputs(9858) <= not(layer0_outputs(8588));
    layer1_outputs(9859) <= (layer0_outputs(765)) xor (layer0_outputs(1684));
    layer1_outputs(9860) <= not(layer0_outputs(7638));
    layer1_outputs(9861) <= not(layer0_outputs(1999));
    layer1_outputs(9862) <= not((layer0_outputs(4531)) and (layer0_outputs(8383)));
    layer1_outputs(9863) <= not((layer0_outputs(6758)) and (layer0_outputs(5261)));
    layer1_outputs(9864) <= not(layer0_outputs(416)) or (layer0_outputs(6159));
    layer1_outputs(9865) <= not(layer0_outputs(1058)) or (layer0_outputs(5765));
    layer1_outputs(9866) <= '0';
    layer1_outputs(9867) <= layer0_outputs(5553);
    layer1_outputs(9868) <= not(layer0_outputs(3777)) or (layer0_outputs(6250));
    layer1_outputs(9869) <= layer0_outputs(3124);
    layer1_outputs(9870) <= (layer0_outputs(3327)) xor (layer0_outputs(474));
    layer1_outputs(9871) <= (layer0_outputs(3801)) or (layer0_outputs(8166));
    layer1_outputs(9872) <= '1';
    layer1_outputs(9873) <= not(layer0_outputs(531));
    layer1_outputs(9874) <= not(layer0_outputs(10217));
    layer1_outputs(9875) <= not(layer0_outputs(1388)) or (layer0_outputs(3995));
    layer1_outputs(9876) <= (layer0_outputs(1220)) and not (layer0_outputs(1383));
    layer1_outputs(9877) <= not((layer0_outputs(4928)) and (layer0_outputs(2160)));
    layer1_outputs(9878) <= (layer0_outputs(2066)) and not (layer0_outputs(727));
    layer1_outputs(9879) <= not((layer0_outputs(2488)) xor (layer0_outputs(2504)));
    layer1_outputs(9880) <= (layer0_outputs(7358)) and not (layer0_outputs(6184));
    layer1_outputs(9881) <= (layer0_outputs(8726)) and not (layer0_outputs(3953));
    layer1_outputs(9882) <= layer0_outputs(4719);
    layer1_outputs(9883) <= layer0_outputs(2210);
    layer1_outputs(9884) <= not(layer0_outputs(9367));
    layer1_outputs(9885) <= (layer0_outputs(1668)) and not (layer0_outputs(2914));
    layer1_outputs(9886) <= '1';
    layer1_outputs(9887) <= layer0_outputs(6166);
    layer1_outputs(9888) <= not(layer0_outputs(9106)) or (layer0_outputs(7963));
    layer1_outputs(9889) <= layer0_outputs(5783);
    layer1_outputs(9890) <= not((layer0_outputs(6706)) and (layer0_outputs(2413)));
    layer1_outputs(9891) <= not((layer0_outputs(1604)) xor (layer0_outputs(6288)));
    layer1_outputs(9892) <= (layer0_outputs(5140)) xor (layer0_outputs(9051));
    layer1_outputs(9893) <= not(layer0_outputs(6814));
    layer1_outputs(9894) <= (layer0_outputs(4287)) and not (layer0_outputs(1244));
    layer1_outputs(9895) <= not(layer0_outputs(9738)) or (layer0_outputs(3122));
    layer1_outputs(9896) <= not((layer0_outputs(2634)) or (layer0_outputs(9836)));
    layer1_outputs(9897) <= (layer0_outputs(5923)) and not (layer0_outputs(8206));
    layer1_outputs(9898) <= layer0_outputs(7619);
    layer1_outputs(9899) <= layer0_outputs(2905);
    layer1_outputs(9900) <= (layer0_outputs(8326)) and not (layer0_outputs(2482));
    layer1_outputs(9901) <= not(layer0_outputs(5630));
    layer1_outputs(9902) <= not(layer0_outputs(6113));
    layer1_outputs(9903) <= (layer0_outputs(7520)) xor (layer0_outputs(1008));
    layer1_outputs(9904) <= not(layer0_outputs(5397)) or (layer0_outputs(118));
    layer1_outputs(9905) <= (layer0_outputs(1920)) and not (layer0_outputs(924));
    layer1_outputs(9906) <= '1';
    layer1_outputs(9907) <= not((layer0_outputs(2791)) xor (layer0_outputs(3711)));
    layer1_outputs(9908) <= not(layer0_outputs(6273));
    layer1_outputs(9909) <= not((layer0_outputs(1147)) and (layer0_outputs(9989)));
    layer1_outputs(9910) <= (layer0_outputs(2661)) and (layer0_outputs(4459));
    layer1_outputs(9911) <= not(layer0_outputs(4035)) or (layer0_outputs(796));
    layer1_outputs(9912) <= not((layer0_outputs(7596)) xor (layer0_outputs(4949)));
    layer1_outputs(9913) <= not((layer0_outputs(8968)) xor (layer0_outputs(4963)));
    layer1_outputs(9914) <= not(layer0_outputs(323));
    layer1_outputs(9915) <= layer0_outputs(7299);
    layer1_outputs(9916) <= not((layer0_outputs(8868)) and (layer0_outputs(1633)));
    layer1_outputs(9917) <= layer0_outputs(2967);
    layer1_outputs(9918) <= '1';
    layer1_outputs(9919) <= layer0_outputs(5623);
    layer1_outputs(9920) <= not((layer0_outputs(664)) and (layer0_outputs(1048)));
    layer1_outputs(9921) <= layer0_outputs(1786);
    layer1_outputs(9922) <= (layer0_outputs(9805)) and not (layer0_outputs(2822));
    layer1_outputs(9923) <= layer0_outputs(8821);
    layer1_outputs(9924) <= not(layer0_outputs(966)) or (layer0_outputs(2037));
    layer1_outputs(9925) <= (layer0_outputs(5815)) and (layer0_outputs(3185));
    layer1_outputs(9926) <= (layer0_outputs(2461)) or (layer0_outputs(8623));
    layer1_outputs(9927) <= not(layer0_outputs(707));
    layer1_outputs(9928) <= '0';
    layer1_outputs(9929) <= '1';
    layer1_outputs(9930) <= (layer0_outputs(3112)) xor (layer0_outputs(4668));
    layer1_outputs(9931) <= not((layer0_outputs(595)) and (layer0_outputs(4396)));
    layer1_outputs(9932) <= (layer0_outputs(869)) or (layer0_outputs(1852));
    layer1_outputs(9933) <= (layer0_outputs(1969)) and not (layer0_outputs(9331));
    layer1_outputs(9934) <= not(layer0_outputs(4579)) or (layer0_outputs(1012));
    layer1_outputs(9935) <= layer0_outputs(4959);
    layer1_outputs(9936) <= '1';
    layer1_outputs(9937) <= (layer0_outputs(2078)) xor (layer0_outputs(1774));
    layer1_outputs(9938) <= not((layer0_outputs(3392)) and (layer0_outputs(2712)));
    layer1_outputs(9939) <= (layer0_outputs(2005)) and (layer0_outputs(4391));
    layer1_outputs(9940) <= (layer0_outputs(5774)) xor (layer0_outputs(6683));
    layer1_outputs(9941) <= layer0_outputs(1036);
    layer1_outputs(9942) <= (layer0_outputs(8220)) and (layer0_outputs(2159));
    layer1_outputs(9943) <= not(layer0_outputs(9441));
    layer1_outputs(9944) <= (layer0_outputs(5960)) xor (layer0_outputs(5914));
    layer1_outputs(9945) <= not((layer0_outputs(7481)) xor (layer0_outputs(6011)));
    layer1_outputs(9946) <= layer0_outputs(3281);
    layer1_outputs(9947) <= layer0_outputs(8892);
    layer1_outputs(9948) <= (layer0_outputs(6614)) and not (layer0_outputs(2785));
    layer1_outputs(9949) <= not((layer0_outputs(2217)) or (layer0_outputs(2284)));
    layer1_outputs(9950) <= (layer0_outputs(9499)) or (layer0_outputs(7950));
    layer1_outputs(9951) <= layer0_outputs(4090);
    layer1_outputs(9952) <= not(layer0_outputs(6304)) or (layer0_outputs(4048));
    layer1_outputs(9953) <= not((layer0_outputs(8976)) and (layer0_outputs(5933)));
    layer1_outputs(9954) <= not(layer0_outputs(9643));
    layer1_outputs(9955) <= not((layer0_outputs(1954)) xor (layer0_outputs(5528)));
    layer1_outputs(9956) <= (layer0_outputs(1567)) and not (layer0_outputs(3188));
    layer1_outputs(9957) <= (layer0_outputs(758)) and not (layer0_outputs(5132));
    layer1_outputs(9958) <= (layer0_outputs(9402)) and not (layer0_outputs(3054));
    layer1_outputs(9959) <= (layer0_outputs(6108)) and not (layer0_outputs(4829));
    layer1_outputs(9960) <= layer0_outputs(2934);
    layer1_outputs(9961) <= (layer0_outputs(8341)) and (layer0_outputs(7764));
    layer1_outputs(9962) <= layer0_outputs(83);
    layer1_outputs(9963) <= '1';
    layer1_outputs(9964) <= not(layer0_outputs(3224)) or (layer0_outputs(4815));
    layer1_outputs(9965) <= not(layer0_outputs(3556));
    layer1_outputs(9966) <= (layer0_outputs(1506)) and (layer0_outputs(96));
    layer1_outputs(9967) <= layer0_outputs(9214);
    layer1_outputs(9968) <= not(layer0_outputs(4672));
    layer1_outputs(9969) <= (layer0_outputs(9050)) and (layer0_outputs(2700));
    layer1_outputs(9970) <= (layer0_outputs(7913)) and not (layer0_outputs(10162));
    layer1_outputs(9971) <= layer0_outputs(7255);
    layer1_outputs(9972) <= layer0_outputs(3446);
    layer1_outputs(9973) <= (layer0_outputs(3421)) and (layer0_outputs(590));
    layer1_outputs(9974) <= '1';
    layer1_outputs(9975) <= (layer0_outputs(8750)) or (layer0_outputs(2760));
    layer1_outputs(9976) <= (layer0_outputs(5915)) or (layer0_outputs(7846));
    layer1_outputs(9977) <= not(layer0_outputs(3111));
    layer1_outputs(9978) <= layer0_outputs(8163);
    layer1_outputs(9979) <= not(layer0_outputs(3741));
    layer1_outputs(9980) <= not((layer0_outputs(4600)) xor (layer0_outputs(7946)));
    layer1_outputs(9981) <= (layer0_outputs(9881)) and not (layer0_outputs(655));
    layer1_outputs(9982) <= (layer0_outputs(9148)) xor (layer0_outputs(265));
    layer1_outputs(9983) <= (layer0_outputs(8926)) and not (layer0_outputs(7678));
    layer1_outputs(9984) <= (layer0_outputs(813)) and (layer0_outputs(3230));
    layer1_outputs(9985) <= not((layer0_outputs(8748)) or (layer0_outputs(6576)));
    layer1_outputs(9986) <= (layer0_outputs(5506)) and (layer0_outputs(6627));
    layer1_outputs(9987) <= (layer0_outputs(8480)) xor (layer0_outputs(6793));
    layer1_outputs(9988) <= (layer0_outputs(7774)) or (layer0_outputs(9964));
    layer1_outputs(9989) <= (layer0_outputs(5977)) xor (layer0_outputs(1136));
    layer1_outputs(9990) <= not((layer0_outputs(4192)) or (layer0_outputs(6545)));
    layer1_outputs(9991) <= not(layer0_outputs(4597));
    layer1_outputs(9992) <= layer0_outputs(4106);
    layer1_outputs(9993) <= (layer0_outputs(129)) and not (layer0_outputs(9610));
    layer1_outputs(9994) <= not(layer0_outputs(5403));
    layer1_outputs(9995) <= (layer0_outputs(163)) and not (layer0_outputs(9957));
    layer1_outputs(9996) <= (layer0_outputs(7814)) or (layer0_outputs(1899));
    layer1_outputs(9997) <= (layer0_outputs(573)) and not (layer0_outputs(3976));
    layer1_outputs(9998) <= layer0_outputs(185);
    layer1_outputs(9999) <= not(layer0_outputs(8085));
    layer1_outputs(10000) <= not(layer0_outputs(2410)) or (layer0_outputs(9570));
    layer1_outputs(10001) <= not((layer0_outputs(4110)) and (layer0_outputs(6973)));
    layer1_outputs(10002) <= (layer0_outputs(3571)) or (layer0_outputs(3317));
    layer1_outputs(10003) <= layer0_outputs(9492);
    layer1_outputs(10004) <= not(layer0_outputs(5313));
    layer1_outputs(10005) <= (layer0_outputs(3049)) xor (layer0_outputs(3487));
    layer1_outputs(10006) <= not(layer0_outputs(1498));
    layer1_outputs(10007) <= (layer0_outputs(2574)) and not (layer0_outputs(7126));
    layer1_outputs(10008) <= not(layer0_outputs(639));
    layer1_outputs(10009) <= layer0_outputs(149);
    layer1_outputs(10010) <= not(layer0_outputs(7720)) or (layer0_outputs(4110));
    layer1_outputs(10011) <= not(layer0_outputs(6831));
    layer1_outputs(10012) <= not(layer0_outputs(7880)) or (layer0_outputs(4191));
    layer1_outputs(10013) <= (layer0_outputs(9927)) and not (layer0_outputs(7974));
    layer1_outputs(10014) <= '0';
    layer1_outputs(10015) <= not(layer0_outputs(260));
    layer1_outputs(10016) <= not(layer0_outputs(3226));
    layer1_outputs(10017) <= layer0_outputs(3676);
    layer1_outputs(10018) <= not(layer0_outputs(2256));
    layer1_outputs(10019) <= not((layer0_outputs(2337)) xor (layer0_outputs(4526)));
    layer1_outputs(10020) <= (layer0_outputs(3737)) and not (layer0_outputs(5734));
    layer1_outputs(10021) <= not(layer0_outputs(2873));
    layer1_outputs(10022) <= not(layer0_outputs(9811)) or (layer0_outputs(9037));
    layer1_outputs(10023) <= not((layer0_outputs(7391)) and (layer0_outputs(6033)));
    layer1_outputs(10024) <= (layer0_outputs(5354)) and (layer0_outputs(2865));
    layer1_outputs(10025) <= layer0_outputs(6816);
    layer1_outputs(10026) <= not(layer0_outputs(4356));
    layer1_outputs(10027) <= layer0_outputs(2558);
    layer1_outputs(10028) <= layer0_outputs(7433);
    layer1_outputs(10029) <= '0';
    layer1_outputs(10030) <= '1';
    layer1_outputs(10031) <= not((layer0_outputs(3761)) and (layer0_outputs(99)));
    layer1_outputs(10032) <= not((layer0_outputs(8009)) xor (layer0_outputs(344)));
    layer1_outputs(10033) <= not((layer0_outputs(4052)) and (layer0_outputs(970)));
    layer1_outputs(10034) <= not(layer0_outputs(3890));
    layer1_outputs(10035) <= (layer0_outputs(10159)) xor (layer0_outputs(7807));
    layer1_outputs(10036) <= not(layer0_outputs(8638));
    layer1_outputs(10037) <= layer0_outputs(1446);
    layer1_outputs(10038) <= not((layer0_outputs(3646)) and (layer0_outputs(5583)));
    layer1_outputs(10039) <= not((layer0_outputs(8861)) and (layer0_outputs(8205)));
    layer1_outputs(10040) <= layer0_outputs(487);
    layer1_outputs(10041) <= (layer0_outputs(252)) and not (layer0_outputs(7591));
    layer1_outputs(10042) <= not(layer0_outputs(4592));
    layer1_outputs(10043) <= (layer0_outputs(1430)) and not (layer0_outputs(3991));
    layer1_outputs(10044) <= (layer0_outputs(4301)) xor (layer0_outputs(3294));
    layer1_outputs(10045) <= not((layer0_outputs(788)) and (layer0_outputs(8697)));
    layer1_outputs(10046) <= (layer0_outputs(1725)) and not (layer0_outputs(6800));
    layer1_outputs(10047) <= not(layer0_outputs(8325)) or (layer0_outputs(7873));
    layer1_outputs(10048) <= (layer0_outputs(9457)) and (layer0_outputs(6925));
    layer1_outputs(10049) <= (layer0_outputs(520)) xor (layer0_outputs(5408));
    layer1_outputs(10050) <= not(layer0_outputs(6083)) or (layer0_outputs(4369));
    layer1_outputs(10051) <= layer0_outputs(9588);
    layer1_outputs(10052) <= layer0_outputs(8187);
    layer1_outputs(10053) <= layer0_outputs(7432);
    layer1_outputs(10054) <= (layer0_outputs(7244)) and not (layer0_outputs(6025));
    layer1_outputs(10055) <= not((layer0_outputs(3903)) xor (layer0_outputs(3383)));
    layer1_outputs(10056) <= '1';
    layer1_outputs(10057) <= not(layer0_outputs(5359)) or (layer0_outputs(8770));
    layer1_outputs(10058) <= (layer0_outputs(967)) and (layer0_outputs(1098));
    layer1_outputs(10059) <= not(layer0_outputs(2238));
    layer1_outputs(10060) <= not((layer0_outputs(1279)) xor (layer0_outputs(3987)));
    layer1_outputs(10061) <= '0';
    layer1_outputs(10062) <= (layer0_outputs(2672)) and not (layer0_outputs(5120));
    layer1_outputs(10063) <= not(layer0_outputs(1824));
    layer1_outputs(10064) <= not(layer0_outputs(875));
    layer1_outputs(10065) <= not((layer0_outputs(9825)) and (layer0_outputs(5073)));
    layer1_outputs(10066) <= not(layer0_outputs(4373));
    layer1_outputs(10067) <= not(layer0_outputs(3164)) or (layer0_outputs(8912));
    layer1_outputs(10068) <= not(layer0_outputs(7135));
    layer1_outputs(10069) <= not(layer0_outputs(9472)) or (layer0_outputs(9704));
    layer1_outputs(10070) <= layer0_outputs(5105);
    layer1_outputs(10071) <= layer0_outputs(429);
    layer1_outputs(10072) <= layer0_outputs(10178);
    layer1_outputs(10073) <= (layer0_outputs(5454)) xor (layer0_outputs(6131));
    layer1_outputs(10074) <= not(layer0_outputs(2749)) or (layer0_outputs(8437));
    layer1_outputs(10075) <= layer0_outputs(3879);
    layer1_outputs(10076) <= not(layer0_outputs(3329)) or (layer0_outputs(1854));
    layer1_outputs(10077) <= not((layer0_outputs(6339)) or (layer0_outputs(2835)));
    layer1_outputs(10078) <= not((layer0_outputs(8815)) or (layer0_outputs(3031)));
    layer1_outputs(10079) <= not(layer0_outputs(9084)) or (layer0_outputs(2805));
    layer1_outputs(10080) <= (layer0_outputs(4344)) or (layer0_outputs(135));
    layer1_outputs(10081) <= layer0_outputs(5964);
    layer1_outputs(10082) <= not(layer0_outputs(5863)) or (layer0_outputs(9756));
    layer1_outputs(10083) <= (layer0_outputs(4361)) or (layer0_outputs(9517));
    layer1_outputs(10084) <= not(layer0_outputs(2947));
    layer1_outputs(10085) <= layer0_outputs(3968);
    layer1_outputs(10086) <= (layer0_outputs(2843)) and not (layer0_outputs(10195));
    layer1_outputs(10087) <= (layer0_outputs(3413)) and (layer0_outputs(6429));
    layer1_outputs(10088) <= not(layer0_outputs(8653));
    layer1_outputs(10089) <= (layer0_outputs(3836)) and not (layer0_outputs(3199));
    layer1_outputs(10090) <= not(layer0_outputs(8123)) or (layer0_outputs(3885));
    layer1_outputs(10091) <= not(layer0_outputs(661));
    layer1_outputs(10092) <= not(layer0_outputs(9551));
    layer1_outputs(10093) <= (layer0_outputs(4913)) and (layer0_outputs(5063));
    layer1_outputs(10094) <= not((layer0_outputs(1543)) or (layer0_outputs(4170)));
    layer1_outputs(10095) <= (layer0_outputs(6129)) xor (layer0_outputs(8402));
    layer1_outputs(10096) <= not(layer0_outputs(1592)) or (layer0_outputs(9074));
    layer1_outputs(10097) <= (layer0_outputs(6361)) and not (layer0_outputs(6970));
    layer1_outputs(10098) <= layer0_outputs(5521);
    layer1_outputs(10099) <= (layer0_outputs(3826)) and (layer0_outputs(9071));
    layer1_outputs(10100) <= not(layer0_outputs(4333)) or (layer0_outputs(8967));
    layer1_outputs(10101) <= layer0_outputs(3333);
    layer1_outputs(10102) <= layer0_outputs(4257);
    layer1_outputs(10103) <= not((layer0_outputs(8026)) or (layer0_outputs(7245)));
    layer1_outputs(10104) <= layer0_outputs(2901);
    layer1_outputs(10105) <= not(layer0_outputs(4058));
    layer1_outputs(10106) <= not(layer0_outputs(9924));
    layer1_outputs(10107) <= not((layer0_outputs(1492)) or (layer0_outputs(3713)));
    layer1_outputs(10108) <= (layer0_outputs(9683)) or (layer0_outputs(6054));
    layer1_outputs(10109) <= (layer0_outputs(5974)) and (layer0_outputs(4504));
    layer1_outputs(10110) <= not(layer0_outputs(7835));
    layer1_outputs(10111) <= layer0_outputs(2443);
    layer1_outputs(10112) <= not(layer0_outputs(4380));
    layer1_outputs(10113) <= (layer0_outputs(2499)) or (layer0_outputs(7487));
    layer1_outputs(10114) <= not(layer0_outputs(3344));
    layer1_outputs(10115) <= (layer0_outputs(9632)) and not (layer0_outputs(5836));
    layer1_outputs(10116) <= '0';
    layer1_outputs(10117) <= (layer0_outputs(3762)) and (layer0_outputs(1972));
    layer1_outputs(10118) <= not(layer0_outputs(3655)) or (layer0_outputs(2069));
    layer1_outputs(10119) <= layer0_outputs(9337);
    layer1_outputs(10120) <= (layer0_outputs(697)) or (layer0_outputs(10092));
    layer1_outputs(10121) <= not(layer0_outputs(7354));
    layer1_outputs(10122) <= layer0_outputs(7486);
    layer1_outputs(10123) <= not(layer0_outputs(4086));
    layer1_outputs(10124) <= layer0_outputs(1278);
    layer1_outputs(10125) <= not(layer0_outputs(8140));
    layer1_outputs(10126) <= not(layer0_outputs(8004));
    layer1_outputs(10127) <= (layer0_outputs(5422)) and not (layer0_outputs(9584));
    layer1_outputs(10128) <= layer0_outputs(751);
    layer1_outputs(10129) <= not((layer0_outputs(9030)) xor (layer0_outputs(951)));
    layer1_outputs(10130) <= (layer0_outputs(6350)) or (layer0_outputs(2144));
    layer1_outputs(10131) <= not(layer0_outputs(539));
    layer1_outputs(10132) <= not(layer0_outputs(7806)) or (layer0_outputs(8137));
    layer1_outputs(10133) <= (layer0_outputs(3165)) and (layer0_outputs(9750));
    layer1_outputs(10134) <= layer0_outputs(7705);
    layer1_outputs(10135) <= (layer0_outputs(7937)) and not (layer0_outputs(7286));
    layer1_outputs(10136) <= (layer0_outputs(9740)) and (layer0_outputs(651));
    layer1_outputs(10137) <= not((layer0_outputs(6402)) or (layer0_outputs(8656)));
    layer1_outputs(10138) <= layer0_outputs(9882);
    layer1_outputs(10139) <= not(layer0_outputs(6234)) or (layer0_outputs(139));
    layer1_outputs(10140) <= layer0_outputs(7143);
    layer1_outputs(10141) <= (layer0_outputs(10217)) and (layer0_outputs(5865));
    layer1_outputs(10142) <= layer0_outputs(1608);
    layer1_outputs(10143) <= (layer0_outputs(4294)) and (layer0_outputs(8648));
    layer1_outputs(10144) <= not(layer0_outputs(188));
    layer1_outputs(10145) <= (layer0_outputs(8337)) or (layer0_outputs(1203));
    layer1_outputs(10146) <= layer0_outputs(4334);
    layer1_outputs(10147) <= not(layer0_outputs(1305));
    layer1_outputs(10148) <= not(layer0_outputs(3149)) or (layer0_outputs(4942));
    layer1_outputs(10149) <= not((layer0_outputs(10091)) and (layer0_outputs(9606)));
    layer1_outputs(10150) <= layer0_outputs(7014);
    layer1_outputs(10151) <= (layer0_outputs(409)) and (layer0_outputs(4366));
    layer1_outputs(10152) <= not(layer0_outputs(7667)) or (layer0_outputs(5809));
    layer1_outputs(10153) <= layer0_outputs(1251);
    layer1_outputs(10154) <= not((layer0_outputs(4337)) xor (layer0_outputs(7664)));
    layer1_outputs(10155) <= not((layer0_outputs(4476)) xor (layer0_outputs(8740)));
    layer1_outputs(10156) <= '1';
    layer1_outputs(10157) <= (layer0_outputs(3637)) xor (layer0_outputs(8864));
    layer1_outputs(10158) <= not((layer0_outputs(6967)) and (layer0_outputs(4412)));
    layer1_outputs(10159) <= not(layer0_outputs(2460));
    layer1_outputs(10160) <= (layer0_outputs(7886)) and not (layer0_outputs(6551));
    layer1_outputs(10161) <= layer0_outputs(71);
    layer1_outputs(10162) <= (layer0_outputs(8247)) or (layer0_outputs(9317));
    layer1_outputs(10163) <= layer0_outputs(6964);
    layer1_outputs(10164) <= layer0_outputs(9915);
    layer1_outputs(10165) <= not(layer0_outputs(5666));
    layer1_outputs(10166) <= (layer0_outputs(7711)) and (layer0_outputs(340));
    layer1_outputs(10167) <= not(layer0_outputs(6438));
    layer1_outputs(10168) <= not(layer0_outputs(8390)) or (layer0_outputs(21));
    layer1_outputs(10169) <= layer0_outputs(9047);
    layer1_outputs(10170) <= layer0_outputs(10215);
    layer1_outputs(10171) <= layer0_outputs(1759);
    layer1_outputs(10172) <= layer0_outputs(5633);
    layer1_outputs(10173) <= not(layer0_outputs(9892));
    layer1_outputs(10174) <= not((layer0_outputs(9974)) and (layer0_outputs(8039)));
    layer1_outputs(10175) <= layer0_outputs(913);
    layer1_outputs(10176) <= (layer0_outputs(2246)) and not (layer0_outputs(9958));
    layer1_outputs(10177) <= not(layer0_outputs(1642)) or (layer0_outputs(789));
    layer1_outputs(10178) <= layer0_outputs(2994);
    layer1_outputs(10179) <= '1';
    layer1_outputs(10180) <= layer0_outputs(4948);
    layer1_outputs(10181) <= not(layer0_outputs(9585));
    layer1_outputs(10182) <= '0';
    layer1_outputs(10183) <= not(layer0_outputs(7130));
    layer1_outputs(10184) <= not((layer0_outputs(3318)) or (layer0_outputs(10212)));
    layer1_outputs(10185) <= not((layer0_outputs(2451)) or (layer0_outputs(1798)));
    layer1_outputs(10186) <= not(layer0_outputs(2372));
    layer1_outputs(10187) <= (layer0_outputs(9364)) and (layer0_outputs(6455));
    layer1_outputs(10188) <= layer0_outputs(5502);
    layer1_outputs(10189) <= layer0_outputs(9698);
    layer1_outputs(10190) <= (layer0_outputs(2689)) and not (layer0_outputs(2862));
    layer1_outputs(10191) <= layer0_outputs(6063);
    layer1_outputs(10192) <= not(layer0_outputs(5336));
    layer1_outputs(10193) <= not((layer0_outputs(3741)) and (layer0_outputs(1429)));
    layer1_outputs(10194) <= not(layer0_outputs(4940));
    layer1_outputs(10195) <= '0';
    layer1_outputs(10196) <= not((layer0_outputs(2079)) and (layer0_outputs(3399)));
    layer1_outputs(10197) <= layer0_outputs(4677);
    layer1_outputs(10198) <= not((layer0_outputs(8958)) xor (layer0_outputs(2095)));
    layer1_outputs(10199) <= not(layer0_outputs(9376));
    layer1_outputs(10200) <= not(layer0_outputs(8663)) or (layer0_outputs(1122));
    layer1_outputs(10201) <= (layer0_outputs(1235)) or (layer0_outputs(8882));
    layer1_outputs(10202) <= not(layer0_outputs(9171));
    layer1_outputs(10203) <= layer0_outputs(2923);
    layer1_outputs(10204) <= (layer0_outputs(8228)) and (layer0_outputs(4301));
    layer1_outputs(10205) <= not(layer0_outputs(2559));
    layer1_outputs(10206) <= layer0_outputs(1771);
    layer1_outputs(10207) <= not(layer0_outputs(5814)) or (layer0_outputs(3765));
    layer1_outputs(10208) <= not((layer0_outputs(4268)) xor (layer0_outputs(2955)));
    layer1_outputs(10209) <= layer0_outputs(2789);
    layer1_outputs(10210) <= not(layer0_outputs(5347));
    layer1_outputs(10211) <= (layer0_outputs(4964)) xor (layer0_outputs(7828));
    layer1_outputs(10212) <= '0';
    layer1_outputs(10213) <= (layer0_outputs(4285)) and not (layer0_outputs(4646));
    layer1_outputs(10214) <= layer0_outputs(5229);
    layer1_outputs(10215) <= not((layer0_outputs(9435)) or (layer0_outputs(3541)));
    layer1_outputs(10216) <= not(layer0_outputs(6090));
    layer1_outputs(10217) <= (layer0_outputs(9653)) and not (layer0_outputs(6981));
    layer1_outputs(10218) <= (layer0_outputs(7934)) and not (layer0_outputs(3647));
    layer1_outputs(10219) <= not((layer0_outputs(2361)) or (layer0_outputs(5486)));
    layer1_outputs(10220) <= not(layer0_outputs(2068));
    layer1_outputs(10221) <= (layer0_outputs(9464)) and not (layer0_outputs(3133));
    layer1_outputs(10222) <= not((layer0_outputs(4014)) xor (layer0_outputs(719)));
    layer1_outputs(10223) <= not(layer0_outputs(10045)) or (layer0_outputs(4801));
    layer1_outputs(10224) <= (layer0_outputs(10184)) and not (layer0_outputs(9444));
    layer1_outputs(10225) <= not((layer0_outputs(6353)) and (layer0_outputs(6449)));
    layer1_outputs(10226) <= (layer0_outputs(7526)) or (layer0_outputs(8965));
    layer1_outputs(10227) <= layer0_outputs(4282);
    layer1_outputs(10228) <= not((layer0_outputs(8731)) and (layer0_outputs(1002)));
    layer1_outputs(10229) <= layer0_outputs(2859);
    layer1_outputs(10230) <= not((layer0_outputs(1814)) or (layer0_outputs(1082)));
    layer1_outputs(10231) <= not(layer0_outputs(5589));
    layer1_outputs(10232) <= (layer0_outputs(6272)) and not (layer0_outputs(5761));
    layer1_outputs(10233) <= not((layer0_outputs(3219)) or (layer0_outputs(5758)));
    layer1_outputs(10234) <= not(layer0_outputs(8966));
    layer1_outputs(10235) <= (layer0_outputs(9453)) or (layer0_outputs(6895));
    layer1_outputs(10236) <= (layer0_outputs(10234)) xor (layer0_outputs(9712));
    layer1_outputs(10237) <= not(layer0_outputs(7224));
    layer1_outputs(10238) <= (layer0_outputs(9805)) and (layer0_outputs(1836));
    layer1_outputs(10239) <= layer0_outputs(7590);
    layer2_outputs(0) <= layer1_outputs(7739);
    layer2_outputs(1) <= not(layer1_outputs(3982));
    layer2_outputs(2) <= (layer1_outputs(7490)) or (layer1_outputs(9789));
    layer2_outputs(3) <= '0';
    layer2_outputs(4) <= not((layer1_outputs(5247)) or (layer1_outputs(8980)));
    layer2_outputs(5) <= not(layer1_outputs(9987));
    layer2_outputs(6) <= not((layer1_outputs(10019)) xor (layer1_outputs(4285)));
    layer2_outputs(7) <= not(layer1_outputs(2958));
    layer2_outputs(8) <= layer1_outputs(6071);
    layer2_outputs(9) <= not(layer1_outputs(8713));
    layer2_outputs(10) <= (layer1_outputs(7802)) and (layer1_outputs(8769));
    layer2_outputs(11) <= layer1_outputs(5061);
    layer2_outputs(12) <= not(layer1_outputs(5915));
    layer2_outputs(13) <= not(layer1_outputs(3636)) or (layer1_outputs(8857));
    layer2_outputs(14) <= (layer1_outputs(5642)) and not (layer1_outputs(8810));
    layer2_outputs(15) <= (layer1_outputs(7171)) or (layer1_outputs(5732));
    layer2_outputs(16) <= not((layer1_outputs(2225)) or (layer1_outputs(9726)));
    layer2_outputs(17) <= not(layer1_outputs(8393));
    layer2_outputs(18) <= not(layer1_outputs(1900));
    layer2_outputs(19) <= not(layer1_outputs(3226));
    layer2_outputs(20) <= (layer1_outputs(4481)) and (layer1_outputs(7084));
    layer2_outputs(21) <= not(layer1_outputs(1339));
    layer2_outputs(22) <= not(layer1_outputs(6856));
    layer2_outputs(23) <= not((layer1_outputs(8255)) xor (layer1_outputs(9823)));
    layer2_outputs(24) <= (layer1_outputs(4718)) and not (layer1_outputs(4139));
    layer2_outputs(25) <= (layer1_outputs(6800)) xor (layer1_outputs(615));
    layer2_outputs(26) <= layer1_outputs(5211);
    layer2_outputs(27) <= not((layer1_outputs(9315)) xor (layer1_outputs(8498)));
    layer2_outputs(28) <= not((layer1_outputs(3008)) or (layer1_outputs(1262)));
    layer2_outputs(29) <= layer1_outputs(845);
    layer2_outputs(30) <= not(layer1_outputs(3879));
    layer2_outputs(31) <= not(layer1_outputs(9206));
    layer2_outputs(32) <= not(layer1_outputs(2554));
    layer2_outputs(33) <= (layer1_outputs(7323)) and (layer1_outputs(7819));
    layer2_outputs(34) <= not(layer1_outputs(2017));
    layer2_outputs(35) <= not((layer1_outputs(3479)) xor (layer1_outputs(5461)));
    layer2_outputs(36) <= not((layer1_outputs(8458)) xor (layer1_outputs(7190)));
    layer2_outputs(37) <= not(layer1_outputs(658));
    layer2_outputs(38) <= not(layer1_outputs(4734));
    layer2_outputs(39) <= not(layer1_outputs(8804));
    layer2_outputs(40) <= not(layer1_outputs(858));
    layer2_outputs(41) <= (layer1_outputs(7961)) xor (layer1_outputs(5209));
    layer2_outputs(42) <= not((layer1_outputs(6441)) and (layer1_outputs(3643)));
    layer2_outputs(43) <= layer1_outputs(27);
    layer2_outputs(44) <= layer1_outputs(8935);
    layer2_outputs(45) <= (layer1_outputs(1442)) and not (layer1_outputs(8151));
    layer2_outputs(46) <= not(layer1_outputs(7558)) or (layer1_outputs(8336));
    layer2_outputs(47) <= not((layer1_outputs(7183)) and (layer1_outputs(2523)));
    layer2_outputs(48) <= not(layer1_outputs(6454));
    layer2_outputs(49) <= not(layer1_outputs(7567)) or (layer1_outputs(1725));
    layer2_outputs(50) <= not(layer1_outputs(1160));
    layer2_outputs(51) <= layer1_outputs(200);
    layer2_outputs(52) <= not(layer1_outputs(2909));
    layer2_outputs(53) <= (layer1_outputs(2826)) or (layer1_outputs(6951));
    layer2_outputs(54) <= (layer1_outputs(1223)) or (layer1_outputs(602));
    layer2_outputs(55) <= (layer1_outputs(1009)) and not (layer1_outputs(8674));
    layer2_outputs(56) <= not((layer1_outputs(9268)) or (layer1_outputs(5399)));
    layer2_outputs(57) <= (layer1_outputs(1442)) and not (layer1_outputs(5067));
    layer2_outputs(58) <= (layer1_outputs(5811)) xor (layer1_outputs(6214));
    layer2_outputs(59) <= (layer1_outputs(788)) or (layer1_outputs(2844));
    layer2_outputs(60) <= layer1_outputs(1249);
    layer2_outputs(61) <= not(layer1_outputs(8154));
    layer2_outputs(62) <= layer1_outputs(3715);
    layer2_outputs(63) <= (layer1_outputs(1315)) or (layer1_outputs(2048));
    layer2_outputs(64) <= (layer1_outputs(10035)) or (layer1_outputs(852));
    layer2_outputs(65) <= not(layer1_outputs(1074));
    layer2_outputs(66) <= layer1_outputs(5816);
    layer2_outputs(67) <= not(layer1_outputs(8968));
    layer2_outputs(68) <= '1';
    layer2_outputs(69) <= not(layer1_outputs(4942));
    layer2_outputs(70) <= (layer1_outputs(6705)) and (layer1_outputs(5589));
    layer2_outputs(71) <= not((layer1_outputs(544)) and (layer1_outputs(1448)));
    layer2_outputs(72) <= (layer1_outputs(3260)) or (layer1_outputs(4056));
    layer2_outputs(73) <= (layer1_outputs(933)) xor (layer1_outputs(5413));
    layer2_outputs(74) <= layer1_outputs(8330);
    layer2_outputs(75) <= not(layer1_outputs(684)) or (layer1_outputs(449));
    layer2_outputs(76) <= layer1_outputs(9831);
    layer2_outputs(77) <= layer1_outputs(4535);
    layer2_outputs(78) <= not(layer1_outputs(9750));
    layer2_outputs(79) <= not((layer1_outputs(7105)) xor (layer1_outputs(8438)));
    layer2_outputs(80) <= not(layer1_outputs(9116));
    layer2_outputs(81) <= (layer1_outputs(9393)) xor (layer1_outputs(4309));
    layer2_outputs(82) <= not((layer1_outputs(1653)) and (layer1_outputs(9824)));
    layer2_outputs(83) <= not(layer1_outputs(3913)) or (layer1_outputs(5210));
    layer2_outputs(84) <= not(layer1_outputs(5503));
    layer2_outputs(85) <= not((layer1_outputs(7664)) xor (layer1_outputs(9412)));
    layer2_outputs(86) <= layer1_outputs(6354);
    layer2_outputs(87) <= layer1_outputs(404);
    layer2_outputs(88) <= not(layer1_outputs(2464)) or (layer1_outputs(7576));
    layer2_outputs(89) <= not(layer1_outputs(1886));
    layer2_outputs(90) <= not((layer1_outputs(8030)) and (layer1_outputs(9325)));
    layer2_outputs(91) <= (layer1_outputs(4552)) and not (layer1_outputs(9611));
    layer2_outputs(92) <= not((layer1_outputs(3714)) and (layer1_outputs(7325)));
    layer2_outputs(93) <= not((layer1_outputs(3049)) xor (layer1_outputs(2370)));
    layer2_outputs(94) <= not((layer1_outputs(7979)) or (layer1_outputs(360)));
    layer2_outputs(95) <= not(layer1_outputs(9087)) or (layer1_outputs(5008));
    layer2_outputs(96) <= not(layer1_outputs(6220)) or (layer1_outputs(8026));
    layer2_outputs(97) <= not(layer1_outputs(4742));
    layer2_outputs(98) <= layer1_outputs(3810);
    layer2_outputs(99) <= not((layer1_outputs(4788)) xor (layer1_outputs(2925)));
    layer2_outputs(100) <= not(layer1_outputs(1461));
    layer2_outputs(101) <= not((layer1_outputs(3524)) xor (layer1_outputs(7441)));
    layer2_outputs(102) <= not(layer1_outputs(2339));
    layer2_outputs(103) <= not(layer1_outputs(1576));
    layer2_outputs(104) <= (layer1_outputs(4522)) and not (layer1_outputs(6290));
    layer2_outputs(105) <= not(layer1_outputs(1187));
    layer2_outputs(106) <= (layer1_outputs(4978)) xor (layer1_outputs(4705));
    layer2_outputs(107) <= (layer1_outputs(4725)) xor (layer1_outputs(5948));
    layer2_outputs(108) <= not((layer1_outputs(1078)) or (layer1_outputs(3619)));
    layer2_outputs(109) <= (layer1_outputs(6918)) xor (layer1_outputs(2965));
    layer2_outputs(110) <= (layer1_outputs(7888)) or (layer1_outputs(2688));
    layer2_outputs(111) <= (layer1_outputs(2951)) and not (layer1_outputs(9808));
    layer2_outputs(112) <= not(layer1_outputs(8504)) or (layer1_outputs(4690));
    layer2_outputs(113) <= layer1_outputs(1357);
    layer2_outputs(114) <= layer1_outputs(4530);
    layer2_outputs(115) <= not(layer1_outputs(613));
    layer2_outputs(116) <= (layer1_outputs(10079)) and not (layer1_outputs(2539));
    layer2_outputs(117) <= layer1_outputs(8693);
    layer2_outputs(118) <= (layer1_outputs(4326)) and (layer1_outputs(3024));
    layer2_outputs(119) <= layer1_outputs(2511);
    layer2_outputs(120) <= (layer1_outputs(3716)) or (layer1_outputs(5043));
    layer2_outputs(121) <= (layer1_outputs(9912)) xor (layer1_outputs(1378));
    layer2_outputs(122) <= not(layer1_outputs(10166)) or (layer1_outputs(7771));
    layer2_outputs(123) <= (layer1_outputs(1766)) or (layer1_outputs(7330));
    layer2_outputs(124) <= not((layer1_outputs(4461)) xor (layer1_outputs(2073)));
    layer2_outputs(125) <= not((layer1_outputs(8358)) and (layer1_outputs(6765)));
    layer2_outputs(126) <= layer1_outputs(7950);
    layer2_outputs(127) <= not(layer1_outputs(6117));
    layer2_outputs(128) <= (layer1_outputs(4642)) and (layer1_outputs(6995));
    layer2_outputs(129) <= layer1_outputs(3300);
    layer2_outputs(130) <= layer1_outputs(8955);
    layer2_outputs(131) <= (layer1_outputs(1890)) and not (layer1_outputs(7669));
    layer2_outputs(132) <= not((layer1_outputs(5279)) or (layer1_outputs(1767)));
    layer2_outputs(133) <= not((layer1_outputs(2967)) or (layer1_outputs(9224)));
    layer2_outputs(134) <= (layer1_outputs(1555)) and not (layer1_outputs(6756));
    layer2_outputs(135) <= layer1_outputs(3120);
    layer2_outputs(136) <= layer1_outputs(9679);
    layer2_outputs(137) <= not((layer1_outputs(5079)) xor (layer1_outputs(8955)));
    layer2_outputs(138) <= not(layer1_outputs(593)) or (layer1_outputs(806));
    layer2_outputs(139) <= not(layer1_outputs(2842)) or (layer1_outputs(6247));
    layer2_outputs(140) <= (layer1_outputs(1356)) and not (layer1_outputs(7443));
    layer2_outputs(141) <= not(layer1_outputs(9910)) or (layer1_outputs(5920));
    layer2_outputs(142) <= not((layer1_outputs(6285)) and (layer1_outputs(6178)));
    layer2_outputs(143) <= layer1_outputs(1003);
    layer2_outputs(144) <= layer1_outputs(9704);
    layer2_outputs(145) <= not(layer1_outputs(6646)) or (layer1_outputs(3458));
    layer2_outputs(146) <= not(layer1_outputs(3092));
    layer2_outputs(147) <= not(layer1_outputs(1488)) or (layer1_outputs(8128));
    layer2_outputs(148) <= not((layer1_outputs(4020)) and (layer1_outputs(4138)));
    layer2_outputs(149) <= (layer1_outputs(712)) and not (layer1_outputs(347));
    layer2_outputs(150) <= layer1_outputs(9505);
    layer2_outputs(151) <= (layer1_outputs(4722)) and (layer1_outputs(8003));
    layer2_outputs(152) <= layer1_outputs(2259);
    layer2_outputs(153) <= not((layer1_outputs(2118)) xor (layer1_outputs(532)));
    layer2_outputs(154) <= (layer1_outputs(420)) and not (layer1_outputs(5038));
    layer2_outputs(155) <= (layer1_outputs(7089)) and not (layer1_outputs(6901));
    layer2_outputs(156) <= (layer1_outputs(6881)) and not (layer1_outputs(9842));
    layer2_outputs(157) <= (layer1_outputs(6220)) or (layer1_outputs(2490));
    layer2_outputs(158) <= layer1_outputs(10051);
    layer2_outputs(159) <= not(layer1_outputs(316));
    layer2_outputs(160) <= layer1_outputs(3901);
    layer2_outputs(161) <= layer1_outputs(10107);
    layer2_outputs(162) <= (layer1_outputs(3927)) xor (layer1_outputs(4784));
    layer2_outputs(163) <= layer1_outputs(3386);
    layer2_outputs(164) <= not((layer1_outputs(139)) or (layer1_outputs(6502)));
    layer2_outputs(165) <= not(layer1_outputs(1006));
    layer2_outputs(166) <= layer1_outputs(9810);
    layer2_outputs(167) <= not((layer1_outputs(8014)) or (layer1_outputs(2407)));
    layer2_outputs(168) <= (layer1_outputs(3224)) and not (layer1_outputs(3387));
    layer2_outputs(169) <= not(layer1_outputs(7747));
    layer2_outputs(170) <= not(layer1_outputs(4081));
    layer2_outputs(171) <= not((layer1_outputs(1439)) or (layer1_outputs(9757)));
    layer2_outputs(172) <= not(layer1_outputs(10000));
    layer2_outputs(173) <= (layer1_outputs(6272)) and (layer1_outputs(4279));
    layer2_outputs(174) <= layer1_outputs(2878);
    layer2_outputs(175) <= not(layer1_outputs(7426));
    layer2_outputs(176) <= not(layer1_outputs(2088));
    layer2_outputs(177) <= (layer1_outputs(882)) or (layer1_outputs(7880));
    layer2_outputs(178) <= layer1_outputs(6509);
    layer2_outputs(179) <= not(layer1_outputs(9242));
    layer2_outputs(180) <= not(layer1_outputs(1971)) or (layer1_outputs(4974));
    layer2_outputs(181) <= not(layer1_outputs(4771));
    layer2_outputs(182) <= not(layer1_outputs(6238));
    layer2_outputs(183) <= layer1_outputs(5503);
    layer2_outputs(184) <= not((layer1_outputs(118)) xor (layer1_outputs(5468)));
    layer2_outputs(185) <= not((layer1_outputs(7996)) and (layer1_outputs(5171)));
    layer2_outputs(186) <= layer1_outputs(187);
    layer2_outputs(187) <= not((layer1_outputs(2064)) or (layer1_outputs(2301)));
    layer2_outputs(188) <= not((layer1_outputs(7478)) xor (layer1_outputs(7033)));
    layer2_outputs(189) <= not(layer1_outputs(7475));
    layer2_outputs(190) <= (layer1_outputs(7389)) and (layer1_outputs(5318));
    layer2_outputs(191) <= layer1_outputs(3625);
    layer2_outputs(192) <= layer1_outputs(10067);
    layer2_outputs(193) <= not(layer1_outputs(96));
    layer2_outputs(194) <= layer1_outputs(5171);
    layer2_outputs(195) <= not(layer1_outputs(2851));
    layer2_outputs(196) <= layer1_outputs(5947);
    layer2_outputs(197) <= not(layer1_outputs(3004));
    layer2_outputs(198) <= not(layer1_outputs(2910));
    layer2_outputs(199) <= layer1_outputs(8137);
    layer2_outputs(200) <= layer1_outputs(942);
    layer2_outputs(201) <= not((layer1_outputs(5252)) or (layer1_outputs(5611)));
    layer2_outputs(202) <= (layer1_outputs(8813)) and (layer1_outputs(4541));
    layer2_outputs(203) <= not(layer1_outputs(4618));
    layer2_outputs(204) <= not(layer1_outputs(2174));
    layer2_outputs(205) <= not(layer1_outputs(3781));
    layer2_outputs(206) <= not(layer1_outputs(6921)) or (layer1_outputs(5861));
    layer2_outputs(207) <= (layer1_outputs(1086)) or (layer1_outputs(4854));
    layer2_outputs(208) <= not(layer1_outputs(9795));
    layer2_outputs(209) <= (layer1_outputs(1048)) xor (layer1_outputs(7346));
    layer2_outputs(210) <= not((layer1_outputs(4779)) xor (layer1_outputs(7403)));
    layer2_outputs(211) <= layer1_outputs(7101);
    layer2_outputs(212) <= (layer1_outputs(4341)) and not (layer1_outputs(1380));
    layer2_outputs(213) <= not(layer1_outputs(7779)) or (layer1_outputs(10087));
    layer2_outputs(214) <= not((layer1_outputs(212)) and (layer1_outputs(4224)));
    layer2_outputs(215) <= (layer1_outputs(4207)) and (layer1_outputs(5720));
    layer2_outputs(216) <= not(layer1_outputs(7430));
    layer2_outputs(217) <= (layer1_outputs(8018)) and not (layer1_outputs(2867));
    layer2_outputs(218) <= not(layer1_outputs(9986));
    layer2_outputs(219) <= layer1_outputs(7122);
    layer2_outputs(220) <= not(layer1_outputs(2740)) or (layer1_outputs(9691));
    layer2_outputs(221) <= (layer1_outputs(9753)) and (layer1_outputs(6352));
    layer2_outputs(222) <= not(layer1_outputs(8973));
    layer2_outputs(223) <= layer1_outputs(5274);
    layer2_outputs(224) <= layer1_outputs(3060);
    layer2_outputs(225) <= '1';
    layer2_outputs(226) <= not((layer1_outputs(7696)) or (layer1_outputs(6972)));
    layer2_outputs(227) <= (layer1_outputs(1812)) or (layer1_outputs(6092));
    layer2_outputs(228) <= not(layer1_outputs(6739));
    layer2_outputs(229) <= layer1_outputs(2463);
    layer2_outputs(230) <= not(layer1_outputs(7642));
    layer2_outputs(231) <= (layer1_outputs(10068)) or (layer1_outputs(5440));
    layer2_outputs(232) <= not(layer1_outputs(1756)) or (layer1_outputs(3896));
    layer2_outputs(233) <= not((layer1_outputs(3524)) xor (layer1_outputs(9250)));
    layer2_outputs(234) <= not(layer1_outputs(1387)) or (layer1_outputs(5684));
    layer2_outputs(235) <= not(layer1_outputs(9323));
    layer2_outputs(236) <= (layer1_outputs(5344)) and not (layer1_outputs(7510));
    layer2_outputs(237) <= (layer1_outputs(3289)) xor (layer1_outputs(3748));
    layer2_outputs(238) <= not(layer1_outputs(6562));
    layer2_outputs(239) <= not(layer1_outputs(4959)) or (layer1_outputs(972));
    layer2_outputs(240) <= (layer1_outputs(5987)) xor (layer1_outputs(6158));
    layer2_outputs(241) <= not((layer1_outputs(8466)) and (layer1_outputs(1205)));
    layer2_outputs(242) <= not(layer1_outputs(4536));
    layer2_outputs(243) <= not(layer1_outputs(2638));
    layer2_outputs(244) <= not(layer1_outputs(1467));
    layer2_outputs(245) <= layer1_outputs(5964);
    layer2_outputs(246) <= not(layer1_outputs(9138));
    layer2_outputs(247) <= not(layer1_outputs(7078));
    layer2_outputs(248) <= (layer1_outputs(5084)) and not (layer1_outputs(7411));
    layer2_outputs(249) <= not(layer1_outputs(79)) or (layer1_outputs(2908));
    layer2_outputs(250) <= not(layer1_outputs(1521));
    layer2_outputs(251) <= layer1_outputs(3114);
    layer2_outputs(252) <= (layer1_outputs(6771)) and not (layer1_outputs(7517));
    layer2_outputs(253) <= not((layer1_outputs(527)) xor (layer1_outputs(9585)));
    layer2_outputs(254) <= not(layer1_outputs(8554));
    layer2_outputs(255) <= layer1_outputs(4540);
    layer2_outputs(256) <= not(layer1_outputs(6690));
    layer2_outputs(257) <= (layer1_outputs(2819)) and (layer1_outputs(8105));
    layer2_outputs(258) <= layer1_outputs(331);
    layer2_outputs(259) <= layer1_outputs(7423);
    layer2_outputs(260) <= not(layer1_outputs(5803));
    layer2_outputs(261) <= layer1_outputs(7851);
    layer2_outputs(262) <= not(layer1_outputs(6558)) or (layer1_outputs(7195));
    layer2_outputs(263) <= (layer1_outputs(881)) or (layer1_outputs(5364));
    layer2_outputs(264) <= layer1_outputs(7515);
    layer2_outputs(265) <= (layer1_outputs(3268)) and not (layer1_outputs(878));
    layer2_outputs(266) <= layer1_outputs(4049);
    layer2_outputs(267) <= not(layer1_outputs(7591));
    layer2_outputs(268) <= (layer1_outputs(3063)) xor (layer1_outputs(9583));
    layer2_outputs(269) <= layer1_outputs(5405);
    layer2_outputs(270) <= not(layer1_outputs(5569)) or (layer1_outputs(6987));
    layer2_outputs(271) <= (layer1_outputs(1383)) and (layer1_outputs(9536));
    layer2_outputs(272) <= layer1_outputs(6317);
    layer2_outputs(273) <= not(layer1_outputs(90));
    layer2_outputs(274) <= layer1_outputs(6245);
    layer2_outputs(275) <= (layer1_outputs(230)) or (layer1_outputs(3876));
    layer2_outputs(276) <= layer1_outputs(5793);
    layer2_outputs(277) <= not(layer1_outputs(5182));
    layer2_outputs(278) <= layer1_outputs(2685);
    layer2_outputs(279) <= not((layer1_outputs(5605)) or (layer1_outputs(8776)));
    layer2_outputs(280) <= not(layer1_outputs(6108)) or (layer1_outputs(8007));
    layer2_outputs(281) <= not(layer1_outputs(2574)) or (layer1_outputs(3557));
    layer2_outputs(282) <= not(layer1_outputs(7831)) or (layer1_outputs(8655));
    layer2_outputs(283) <= (layer1_outputs(6464)) and not (layer1_outputs(4364));
    layer2_outputs(284) <= not((layer1_outputs(2961)) and (layer1_outputs(8784)));
    layer2_outputs(285) <= not(layer1_outputs(454));
    layer2_outputs(286) <= not(layer1_outputs(10107));
    layer2_outputs(287) <= '0';
    layer2_outputs(288) <= not((layer1_outputs(1378)) and (layer1_outputs(4046)));
    layer2_outputs(289) <= (layer1_outputs(4472)) xor (layer1_outputs(3882));
    layer2_outputs(290) <= not(layer1_outputs(9553)) or (layer1_outputs(5088));
    layer2_outputs(291) <= '0';
    layer2_outputs(292) <= layer1_outputs(6794);
    layer2_outputs(293) <= not(layer1_outputs(4856));
    layer2_outputs(294) <= not((layer1_outputs(9665)) or (layer1_outputs(5925)));
    layer2_outputs(295) <= not(layer1_outputs(5345));
    layer2_outputs(296) <= not(layer1_outputs(3072));
    layer2_outputs(297) <= (layer1_outputs(649)) or (layer1_outputs(6462));
    layer2_outputs(298) <= layer1_outputs(8355);
    layer2_outputs(299) <= layer1_outputs(7670);
    layer2_outputs(300) <= layer1_outputs(924);
    layer2_outputs(301) <= not(layer1_outputs(5790));
    layer2_outputs(302) <= not(layer1_outputs(4425));
    layer2_outputs(303) <= (layer1_outputs(7932)) and not (layer1_outputs(1732));
    layer2_outputs(304) <= (layer1_outputs(6554)) and not (layer1_outputs(2764));
    layer2_outputs(305) <= (layer1_outputs(4999)) or (layer1_outputs(1688));
    layer2_outputs(306) <= (layer1_outputs(1336)) and (layer1_outputs(343));
    layer2_outputs(307) <= not(layer1_outputs(2028)) or (layer1_outputs(2893));
    layer2_outputs(308) <= not(layer1_outputs(6725));
    layer2_outputs(309) <= not(layer1_outputs(3428));
    layer2_outputs(310) <= (layer1_outputs(1380)) xor (layer1_outputs(6080));
    layer2_outputs(311) <= (layer1_outputs(9464)) and (layer1_outputs(4658));
    layer2_outputs(312) <= not(layer1_outputs(7737));
    layer2_outputs(313) <= (layer1_outputs(1698)) xor (layer1_outputs(7943));
    layer2_outputs(314) <= not(layer1_outputs(6378)) or (layer1_outputs(5863));
    layer2_outputs(315) <= (layer1_outputs(7118)) xor (layer1_outputs(5263));
    layer2_outputs(316) <= not(layer1_outputs(6957));
    layer2_outputs(317) <= (layer1_outputs(8880)) xor (layer1_outputs(4054));
    layer2_outputs(318) <= (layer1_outputs(7111)) xor (layer1_outputs(3941));
    layer2_outputs(319) <= (layer1_outputs(4026)) and (layer1_outputs(1529));
    layer2_outputs(320) <= (layer1_outputs(3383)) and not (layer1_outputs(806));
    layer2_outputs(321) <= not(layer1_outputs(1811));
    layer2_outputs(322) <= layer1_outputs(1335);
    layer2_outputs(323) <= not(layer1_outputs(9357)) or (layer1_outputs(822));
    layer2_outputs(324) <= (layer1_outputs(7447)) and not (layer1_outputs(4000));
    layer2_outputs(325) <= (layer1_outputs(6786)) and not (layer1_outputs(6943));
    layer2_outputs(326) <= not((layer1_outputs(5996)) xor (layer1_outputs(5263)));
    layer2_outputs(327) <= not(layer1_outputs(1349));
    layer2_outputs(328) <= not((layer1_outputs(4997)) or (layer1_outputs(6194)));
    layer2_outputs(329) <= layer1_outputs(2549);
    layer2_outputs(330) <= layer1_outputs(1450);
    layer2_outputs(331) <= not((layer1_outputs(1341)) and (layer1_outputs(1045)));
    layer2_outputs(332) <= not(layer1_outputs(7238));
    layer2_outputs(333) <= (layer1_outputs(10066)) xor (layer1_outputs(8724));
    layer2_outputs(334) <= not(layer1_outputs(8209)) or (layer1_outputs(555));
    layer2_outputs(335) <= layer1_outputs(8045);
    layer2_outputs(336) <= layer1_outputs(5454);
    layer2_outputs(337) <= (layer1_outputs(7803)) xor (layer1_outputs(3102));
    layer2_outputs(338) <= (layer1_outputs(5086)) and (layer1_outputs(4438));
    layer2_outputs(339) <= not(layer1_outputs(2085));
    layer2_outputs(340) <= not((layer1_outputs(5208)) xor (layer1_outputs(4146)));
    layer2_outputs(341) <= layer1_outputs(646);
    layer2_outputs(342) <= layer1_outputs(428);
    layer2_outputs(343) <= not(layer1_outputs(8990));
    layer2_outputs(344) <= (layer1_outputs(6627)) xor (layer1_outputs(5483));
    layer2_outputs(345) <= (layer1_outputs(3648)) and (layer1_outputs(9332));
    layer2_outputs(346) <= not(layer1_outputs(2572));
    layer2_outputs(347) <= (layer1_outputs(8553)) and not (layer1_outputs(5058));
    layer2_outputs(348) <= not(layer1_outputs(6731));
    layer2_outputs(349) <= not(layer1_outputs(8212));
    layer2_outputs(350) <= (layer1_outputs(8963)) or (layer1_outputs(8678));
    layer2_outputs(351) <= (layer1_outputs(6631)) or (layer1_outputs(1063));
    layer2_outputs(352) <= not((layer1_outputs(4358)) xor (layer1_outputs(7131)));
    layer2_outputs(353) <= not(layer1_outputs(2377));
    layer2_outputs(354) <= not(layer1_outputs(6812));
    layer2_outputs(355) <= not(layer1_outputs(9843));
    layer2_outputs(356) <= not(layer1_outputs(2296));
    layer2_outputs(357) <= layer1_outputs(5908);
    layer2_outputs(358) <= layer1_outputs(9361);
    layer2_outputs(359) <= not(layer1_outputs(9489));
    layer2_outputs(360) <= layer1_outputs(7645);
    layer2_outputs(361) <= not(layer1_outputs(2638));
    layer2_outputs(362) <= not(layer1_outputs(2345));
    layer2_outputs(363) <= not((layer1_outputs(1371)) xor (layer1_outputs(7844)));
    layer2_outputs(364) <= not(layer1_outputs(1176));
    layer2_outputs(365) <= not(layer1_outputs(9656));
    layer2_outputs(366) <= not(layer1_outputs(5789));
    layer2_outputs(367) <= not(layer1_outputs(4195));
    layer2_outputs(368) <= (layer1_outputs(9114)) xor (layer1_outputs(3579));
    layer2_outputs(369) <= not(layer1_outputs(810));
    layer2_outputs(370) <= layer1_outputs(9449);
    layer2_outputs(371) <= layer1_outputs(7524);
    layer2_outputs(372) <= (layer1_outputs(2044)) xor (layer1_outputs(5909));
    layer2_outputs(373) <= (layer1_outputs(6246)) or (layer1_outputs(7695));
    layer2_outputs(374) <= not((layer1_outputs(4439)) or (layer1_outputs(4874)));
    layer2_outputs(375) <= not(layer1_outputs(5989));
    layer2_outputs(376) <= not(layer1_outputs(4565));
    layer2_outputs(377) <= (layer1_outputs(2526)) and not (layer1_outputs(1969));
    layer2_outputs(378) <= not(layer1_outputs(9407));
    layer2_outputs(379) <= (layer1_outputs(2538)) xor (layer1_outputs(4795));
    layer2_outputs(380) <= (layer1_outputs(2922)) xor (layer1_outputs(9442));
    layer2_outputs(381) <= not(layer1_outputs(7070));
    layer2_outputs(382) <= not(layer1_outputs(6336)) or (layer1_outputs(5092));
    layer2_outputs(383) <= not((layer1_outputs(7348)) or (layer1_outputs(3652)));
    layer2_outputs(384) <= '0';
    layer2_outputs(385) <= layer1_outputs(8118);
    layer2_outputs(386) <= (layer1_outputs(1001)) and not (layer1_outputs(9122));
    layer2_outputs(387) <= not((layer1_outputs(3282)) xor (layer1_outputs(3001)));
    layer2_outputs(388) <= layer1_outputs(970);
    layer2_outputs(389) <= (layer1_outputs(1228)) xor (layer1_outputs(6463));
    layer2_outputs(390) <= not((layer1_outputs(10016)) or (layer1_outputs(7748)));
    layer2_outputs(391) <= not(layer1_outputs(7265)) or (layer1_outputs(6672));
    layer2_outputs(392) <= (layer1_outputs(2148)) and not (layer1_outputs(9743));
    layer2_outputs(393) <= layer1_outputs(9643);
    layer2_outputs(394) <= layer1_outputs(3031);
    layer2_outputs(395) <= not(layer1_outputs(8765));
    layer2_outputs(396) <= not(layer1_outputs(1365)) or (layer1_outputs(4043));
    layer2_outputs(397) <= not(layer1_outputs(6478)) or (layer1_outputs(8349));
    layer2_outputs(398) <= (layer1_outputs(6823)) and not (layer1_outputs(3198));
    layer2_outputs(399) <= not((layer1_outputs(4783)) xor (layer1_outputs(7304)));
    layer2_outputs(400) <= not((layer1_outputs(8200)) or (layer1_outputs(8325)));
    layer2_outputs(401) <= layer1_outputs(3798);
    layer2_outputs(402) <= '1';
    layer2_outputs(403) <= not((layer1_outputs(1427)) and (layer1_outputs(9053)));
    layer2_outputs(404) <= layer1_outputs(7228);
    layer2_outputs(405) <= not((layer1_outputs(6596)) or (layer1_outputs(8252)));
    layer2_outputs(406) <= (layer1_outputs(3144)) and not (layer1_outputs(8224));
    layer2_outputs(407) <= (layer1_outputs(5235)) and not (layer1_outputs(5135));
    layer2_outputs(408) <= not(layer1_outputs(6880)) or (layer1_outputs(3907));
    layer2_outputs(409) <= not(layer1_outputs(5945));
    layer2_outputs(410) <= layer1_outputs(3189);
    layer2_outputs(411) <= not((layer1_outputs(4010)) xor (layer1_outputs(5064)));
    layer2_outputs(412) <= layer1_outputs(9767);
    layer2_outputs(413) <= not(layer1_outputs(954));
    layer2_outputs(414) <= layer1_outputs(7186);
    layer2_outputs(415) <= not(layer1_outputs(3829));
    layer2_outputs(416) <= layer1_outputs(3551);
    layer2_outputs(417) <= not((layer1_outputs(4386)) or (layer1_outputs(5231)));
    layer2_outputs(418) <= layer1_outputs(7374);
    layer2_outputs(419) <= layer1_outputs(8073);
    layer2_outputs(420) <= (layer1_outputs(3549)) or (layer1_outputs(7455));
    layer2_outputs(421) <= layer1_outputs(9323);
    layer2_outputs(422) <= layer1_outputs(2774);
    layer2_outputs(423) <= not(layer1_outputs(9676));
    layer2_outputs(424) <= not(layer1_outputs(6162));
    layer2_outputs(425) <= not(layer1_outputs(7747));
    layer2_outputs(426) <= (layer1_outputs(7684)) and not (layer1_outputs(5379));
    layer2_outputs(427) <= not(layer1_outputs(6159));
    layer2_outputs(428) <= not(layer1_outputs(3243));
    layer2_outputs(429) <= not(layer1_outputs(4256));
    layer2_outputs(430) <= not(layer1_outputs(8416)) or (layer1_outputs(9960));
    layer2_outputs(431) <= (layer1_outputs(2758)) and (layer1_outputs(688));
    layer2_outputs(432) <= not((layer1_outputs(7364)) and (layer1_outputs(8014)));
    layer2_outputs(433) <= (layer1_outputs(9432)) or (layer1_outputs(6574));
    layer2_outputs(434) <= not(layer1_outputs(3663)) or (layer1_outputs(8375));
    layer2_outputs(435) <= (layer1_outputs(385)) or (layer1_outputs(9541));
    layer2_outputs(436) <= not(layer1_outputs(298)) or (layer1_outputs(5735));
    layer2_outputs(437) <= layer1_outputs(5961);
    layer2_outputs(438) <= not(layer1_outputs(5224)) or (layer1_outputs(209));
    layer2_outputs(439) <= layer1_outputs(2992);
    layer2_outputs(440) <= not((layer1_outputs(9087)) xor (layer1_outputs(9851)));
    layer2_outputs(441) <= not(layer1_outputs(7561));
    layer2_outputs(442) <= not(layer1_outputs(7871));
    layer2_outputs(443) <= not(layer1_outputs(7476));
    layer2_outputs(444) <= not((layer1_outputs(1352)) xor (layer1_outputs(112)));
    layer2_outputs(445) <= (layer1_outputs(9042)) and not (layer1_outputs(497));
    layer2_outputs(446) <= layer1_outputs(6642);
    layer2_outputs(447) <= layer1_outputs(7299);
    layer2_outputs(448) <= layer1_outputs(890);
    layer2_outputs(449) <= layer1_outputs(6993);
    layer2_outputs(450) <= (layer1_outputs(593)) xor (layer1_outputs(6819));
    layer2_outputs(451) <= layer1_outputs(3017);
    layer2_outputs(452) <= layer1_outputs(4986);
    layer2_outputs(453) <= not(layer1_outputs(3419));
    layer2_outputs(454) <= not(layer1_outputs(4545));
    layer2_outputs(455) <= layer1_outputs(6533);
    layer2_outputs(456) <= not(layer1_outputs(301));
    layer2_outputs(457) <= (layer1_outputs(1698)) and (layer1_outputs(3806));
    layer2_outputs(458) <= (layer1_outputs(6620)) and not (layer1_outputs(4083));
    layer2_outputs(459) <= (layer1_outputs(9722)) and not (layer1_outputs(6757));
    layer2_outputs(460) <= (layer1_outputs(9173)) and (layer1_outputs(8852));
    layer2_outputs(461) <= not(layer1_outputs(8063)) or (layer1_outputs(9370));
    layer2_outputs(462) <= not(layer1_outputs(2419));
    layer2_outputs(463) <= layer1_outputs(1135);
    layer2_outputs(464) <= layer1_outputs(5584);
    layer2_outputs(465) <= not((layer1_outputs(3420)) xor (layer1_outputs(5)));
    layer2_outputs(466) <= not(layer1_outputs(8431));
    layer2_outputs(467) <= not(layer1_outputs(814));
    layer2_outputs(468) <= (layer1_outputs(5623)) and not (layer1_outputs(4960));
    layer2_outputs(469) <= not((layer1_outputs(9184)) and (layer1_outputs(6404)));
    layer2_outputs(470) <= not(layer1_outputs(9953)) or (layer1_outputs(1273));
    layer2_outputs(471) <= not(layer1_outputs(7858)) or (layer1_outputs(7772));
    layer2_outputs(472) <= not(layer1_outputs(4733));
    layer2_outputs(473) <= not(layer1_outputs(9492));
    layer2_outputs(474) <= layer1_outputs(7654);
    layer2_outputs(475) <= (layer1_outputs(5119)) xor (layer1_outputs(2968));
    layer2_outputs(476) <= not((layer1_outputs(3767)) xor (layer1_outputs(3854)));
    layer2_outputs(477) <= not(layer1_outputs(7352));
    layer2_outputs(478) <= layer1_outputs(1334);
    layer2_outputs(479) <= not(layer1_outputs(5496)) or (layer1_outputs(3540));
    layer2_outputs(480) <= layer1_outputs(4316);
    layer2_outputs(481) <= not((layer1_outputs(3506)) and (layer1_outputs(10125)));
    layer2_outputs(482) <= layer1_outputs(594);
    layer2_outputs(483) <= not(layer1_outputs(9923));
    layer2_outputs(484) <= not(layer1_outputs(7461));
    layer2_outputs(485) <= (layer1_outputs(1840)) and not (layer1_outputs(3611));
    layer2_outputs(486) <= not((layer1_outputs(6313)) xor (layer1_outputs(4570)));
    layer2_outputs(487) <= not(layer1_outputs(437));
    layer2_outputs(488) <= (layer1_outputs(1437)) and not (layer1_outputs(1918));
    layer2_outputs(489) <= not(layer1_outputs(8711));
    layer2_outputs(490) <= (layer1_outputs(4417)) and not (layer1_outputs(1183));
    layer2_outputs(491) <= not(layer1_outputs(7171)) or (layer1_outputs(7275));
    layer2_outputs(492) <= not(layer1_outputs(8456));
    layer2_outputs(493) <= not((layer1_outputs(5416)) or (layer1_outputs(2570)));
    layer2_outputs(494) <= layer1_outputs(8918);
    layer2_outputs(495) <= layer1_outputs(4615);
    layer2_outputs(496) <= not((layer1_outputs(1393)) or (layer1_outputs(4840)));
    layer2_outputs(497) <= not(layer1_outputs(293));
    layer2_outputs(498) <= (layer1_outputs(812)) or (layer1_outputs(9305));
    layer2_outputs(499) <= (layer1_outputs(5096)) and not (layer1_outputs(995));
    layer2_outputs(500) <= not(layer1_outputs(7769));
    layer2_outputs(501) <= not((layer1_outputs(112)) xor (layer1_outputs(8600)));
    layer2_outputs(502) <= not((layer1_outputs(3690)) xor (layer1_outputs(1455)));
    layer2_outputs(503) <= not((layer1_outputs(3408)) xor (layer1_outputs(3515)));
    layer2_outputs(504) <= layer1_outputs(1710);
    layer2_outputs(505) <= not(layer1_outputs(4362)) or (layer1_outputs(3534));
    layer2_outputs(506) <= not(layer1_outputs(1392));
    layer2_outputs(507) <= not((layer1_outputs(4828)) xor (layer1_outputs(6307)));
    layer2_outputs(508) <= (layer1_outputs(540)) or (layer1_outputs(1984));
    layer2_outputs(509) <= not(layer1_outputs(7113));
    layer2_outputs(510) <= (layer1_outputs(4001)) and (layer1_outputs(8614));
    layer2_outputs(511) <= layer1_outputs(7151);
    layer2_outputs(512) <= not(layer1_outputs(7066));
    layer2_outputs(513) <= not(layer1_outputs(5697));
    layer2_outputs(514) <= layer1_outputs(2503);
    layer2_outputs(515) <= not(layer1_outputs(9398));
    layer2_outputs(516) <= (layer1_outputs(5913)) and not (layer1_outputs(6375));
    layer2_outputs(517) <= not(layer1_outputs(4791));
    layer2_outputs(518) <= not(layer1_outputs(8520));
    layer2_outputs(519) <= not((layer1_outputs(5251)) xor (layer1_outputs(3050)));
    layer2_outputs(520) <= (layer1_outputs(6763)) xor (layer1_outputs(1645));
    layer2_outputs(521) <= layer1_outputs(7500);
    layer2_outputs(522) <= layer1_outputs(9058);
    layer2_outputs(523) <= not((layer1_outputs(1016)) and (layer1_outputs(790)));
    layer2_outputs(524) <= not((layer1_outputs(2849)) or (layer1_outputs(954)));
    layer2_outputs(525) <= '1';
    layer2_outputs(526) <= (layer1_outputs(2058)) and not (layer1_outputs(579));
    layer2_outputs(527) <= not(layer1_outputs(1935)) or (layer1_outputs(3846));
    layer2_outputs(528) <= not((layer1_outputs(445)) xor (layer1_outputs(2602)));
    layer2_outputs(529) <= layer1_outputs(125);
    layer2_outputs(530) <= not(layer1_outputs(8002)) or (layer1_outputs(2401));
    layer2_outputs(531) <= layer1_outputs(3051);
    layer2_outputs(532) <= (layer1_outputs(4674)) or (layer1_outputs(3755));
    layer2_outputs(533) <= not(layer1_outputs(8116));
    layer2_outputs(534) <= layer1_outputs(1621);
    layer2_outputs(535) <= not((layer1_outputs(6166)) xor (layer1_outputs(6434)));
    layer2_outputs(536) <= not(layer1_outputs(2483));
    layer2_outputs(537) <= (layer1_outputs(8251)) xor (layer1_outputs(9543));
    layer2_outputs(538) <= (layer1_outputs(5565)) and not (layer1_outputs(6041));
    layer2_outputs(539) <= not(layer1_outputs(4332));
    layer2_outputs(540) <= (layer1_outputs(7857)) xor (layer1_outputs(6592));
    layer2_outputs(541) <= layer1_outputs(8922);
    layer2_outputs(542) <= not(layer1_outputs(741));
    layer2_outputs(543) <= (layer1_outputs(4509)) and not (layer1_outputs(2311));
    layer2_outputs(544) <= layer1_outputs(1821);
    layer2_outputs(545) <= not(layer1_outputs(1665)) or (layer1_outputs(1551));
    layer2_outputs(546) <= (layer1_outputs(3033)) xor (layer1_outputs(7101));
    layer2_outputs(547) <= not(layer1_outputs(5422));
    layer2_outputs(548) <= layer1_outputs(4621);
    layer2_outputs(549) <= (layer1_outputs(1049)) and not (layer1_outputs(1867));
    layer2_outputs(550) <= not(layer1_outputs(7974));
    layer2_outputs(551) <= not(layer1_outputs(935));
    layer2_outputs(552) <= layer1_outputs(2851);
    layer2_outputs(553) <= layer1_outputs(6116);
    layer2_outputs(554) <= layer1_outputs(3112);
    layer2_outputs(555) <= not(layer1_outputs(10167));
    layer2_outputs(556) <= layer1_outputs(9830);
    layer2_outputs(557) <= not((layer1_outputs(6497)) xor (layer1_outputs(852)));
    layer2_outputs(558) <= not(layer1_outputs(9511)) or (layer1_outputs(1800));
    layer2_outputs(559) <= not(layer1_outputs(5726));
    layer2_outputs(560) <= not(layer1_outputs(1489));
    layer2_outputs(561) <= not(layer1_outputs(2596));
    layer2_outputs(562) <= not((layer1_outputs(10026)) or (layer1_outputs(3442)));
    layer2_outputs(563) <= not(layer1_outputs(2230));
    layer2_outputs(564) <= layer1_outputs(6085);
    layer2_outputs(565) <= not(layer1_outputs(1429)) or (layer1_outputs(5449));
    layer2_outputs(566) <= (layer1_outputs(10138)) xor (layer1_outputs(2033));
    layer2_outputs(567) <= not((layer1_outputs(6019)) and (layer1_outputs(8624)));
    layer2_outputs(568) <= not(layer1_outputs(2594));
    layer2_outputs(569) <= layer1_outputs(3884);
    layer2_outputs(570) <= not(layer1_outputs(1290)) or (layer1_outputs(3533));
    layer2_outputs(571) <= '1';
    layer2_outputs(572) <= not(layer1_outputs(2433));
    layer2_outputs(573) <= (layer1_outputs(6370)) and not (layer1_outputs(3432));
    layer2_outputs(574) <= not((layer1_outputs(5020)) or (layer1_outputs(4858)));
    layer2_outputs(575) <= layer1_outputs(242);
    layer2_outputs(576) <= (layer1_outputs(7824)) xor (layer1_outputs(8689));
    layer2_outputs(577) <= (layer1_outputs(6594)) or (layer1_outputs(10197));
    layer2_outputs(578) <= (layer1_outputs(5043)) xor (layer1_outputs(1751));
    layer2_outputs(579) <= '1';
    layer2_outputs(580) <= (layer1_outputs(107)) and (layer1_outputs(7266));
    layer2_outputs(581) <= (layer1_outputs(3406)) xor (layer1_outputs(2871));
    layer2_outputs(582) <= layer1_outputs(4446);
    layer2_outputs(583) <= (layer1_outputs(9085)) and not (layer1_outputs(616));
    layer2_outputs(584) <= not((layer1_outputs(3054)) or (layer1_outputs(5697)));
    layer2_outputs(585) <= layer1_outputs(1988);
    layer2_outputs(586) <= not((layer1_outputs(4468)) xor (layer1_outputs(6784)));
    layer2_outputs(587) <= not(layer1_outputs(1668));
    layer2_outputs(588) <= not(layer1_outputs(3790));
    layer2_outputs(589) <= not((layer1_outputs(4296)) xor (layer1_outputs(4022)));
    layer2_outputs(590) <= layer1_outputs(3558);
    layer2_outputs(591) <= (layer1_outputs(10119)) xor (layer1_outputs(9373));
    layer2_outputs(592) <= layer1_outputs(3683);
    layer2_outputs(593) <= not((layer1_outputs(7408)) or (layer1_outputs(7501)));
    layer2_outputs(594) <= not((layer1_outputs(2218)) xor (layer1_outputs(5633)));
    layer2_outputs(595) <= layer1_outputs(10011);
    layer2_outputs(596) <= layer1_outputs(5205);
    layer2_outputs(597) <= layer1_outputs(2043);
    layer2_outputs(598) <= layer1_outputs(2754);
    layer2_outputs(599) <= layer1_outputs(6869);
    layer2_outputs(600) <= not(layer1_outputs(4306));
    layer2_outputs(601) <= not((layer1_outputs(871)) or (layer1_outputs(5771)));
    layer2_outputs(602) <= (layer1_outputs(7874)) xor (layer1_outputs(1611));
    layer2_outputs(603) <= layer1_outputs(32);
    layer2_outputs(604) <= (layer1_outputs(5883)) and not (layer1_outputs(9818));
    layer2_outputs(605) <= layer1_outputs(8174);
    layer2_outputs(606) <= not(layer1_outputs(4229));
    layer2_outputs(607) <= not(layer1_outputs(2785));
    layer2_outputs(608) <= not(layer1_outputs(9816));
    layer2_outputs(609) <= not(layer1_outputs(1871)) or (layer1_outputs(14));
    layer2_outputs(610) <= (layer1_outputs(1596)) xor (layer1_outputs(2938));
    layer2_outputs(611) <= not(layer1_outputs(2834));
    layer2_outputs(612) <= layer1_outputs(1694);
    layer2_outputs(613) <= not(layer1_outputs(2846));
    layer2_outputs(614) <= not(layer1_outputs(1465));
    layer2_outputs(615) <= (layer1_outputs(3564)) xor (layer1_outputs(6569));
    layer2_outputs(616) <= not(layer1_outputs(9706)) or (layer1_outputs(5036));
    layer2_outputs(617) <= layer1_outputs(6562);
    layer2_outputs(618) <= not((layer1_outputs(6397)) xor (layer1_outputs(2388)));
    layer2_outputs(619) <= layer1_outputs(8526);
    layer2_outputs(620) <= layer1_outputs(5719);
    layer2_outputs(621) <= '1';
    layer2_outputs(622) <= layer1_outputs(3572);
    layer2_outputs(623) <= layer1_outputs(621);
    layer2_outputs(624) <= '0';
    layer2_outputs(625) <= not(layer1_outputs(8024)) or (layer1_outputs(4630));
    layer2_outputs(626) <= not(layer1_outputs(6875)) or (layer1_outputs(8411));
    layer2_outputs(627) <= not((layer1_outputs(7392)) or (layer1_outputs(4213)));
    layer2_outputs(628) <= (layer1_outputs(4493)) and not (layer1_outputs(88));
    layer2_outputs(629) <= not((layer1_outputs(441)) or (layer1_outputs(9600)));
    layer2_outputs(630) <= not(layer1_outputs(1333));
    layer2_outputs(631) <= (layer1_outputs(9032)) xor (layer1_outputs(5342));
    layer2_outputs(632) <= not(layer1_outputs(4903));
    layer2_outputs(633) <= (layer1_outputs(7081)) and not (layer1_outputs(8760));
    layer2_outputs(634) <= (layer1_outputs(6044)) and not (layer1_outputs(4100));
    layer2_outputs(635) <= layer1_outputs(8721);
    layer2_outputs(636) <= (layer1_outputs(4538)) and (layer1_outputs(4433));
    layer2_outputs(637) <= not(layer1_outputs(2114));
    layer2_outputs(638) <= layer1_outputs(8718);
    layer2_outputs(639) <= (layer1_outputs(4931)) and not (layer1_outputs(4485));
    layer2_outputs(640) <= (layer1_outputs(7572)) or (layer1_outputs(5094));
    layer2_outputs(641) <= (layer1_outputs(4955)) and not (layer1_outputs(7332));
    layer2_outputs(642) <= not((layer1_outputs(8092)) or (layer1_outputs(10159)));
    layer2_outputs(643) <= layer1_outputs(9507);
    layer2_outputs(644) <= (layer1_outputs(160)) or (layer1_outputs(4612));
    layer2_outputs(645) <= not(layer1_outputs(9799));
    layer2_outputs(646) <= (layer1_outputs(4850)) xor (layer1_outputs(2380));
    layer2_outputs(647) <= layer1_outputs(121);
    layer2_outputs(648) <= (layer1_outputs(6025)) and not (layer1_outputs(1282));
    layer2_outputs(649) <= not((layer1_outputs(121)) xor (layer1_outputs(8916)));
    layer2_outputs(650) <= layer1_outputs(18);
    layer2_outputs(651) <= not(layer1_outputs(9217));
    layer2_outputs(652) <= layer1_outputs(8830);
    layer2_outputs(653) <= not(layer1_outputs(7897));
    layer2_outputs(654) <= not(layer1_outputs(7755));
    layer2_outputs(655) <= not(layer1_outputs(7282));
    layer2_outputs(656) <= not(layer1_outputs(2885));
    layer2_outputs(657) <= (layer1_outputs(6495)) or (layer1_outputs(1848));
    layer2_outputs(658) <= not((layer1_outputs(4183)) xor (layer1_outputs(4709)));
    layer2_outputs(659) <= not((layer1_outputs(2775)) or (layer1_outputs(2792)));
    layer2_outputs(660) <= not((layer1_outputs(2424)) and (layer1_outputs(1688)));
    layer2_outputs(661) <= not(layer1_outputs(2197)) or (layer1_outputs(3130));
    layer2_outputs(662) <= not(layer1_outputs(5190));
    layer2_outputs(663) <= (layer1_outputs(7535)) or (layer1_outputs(8032));
    layer2_outputs(664) <= not((layer1_outputs(1446)) or (layer1_outputs(6182)));
    layer2_outputs(665) <= not(layer1_outputs(1448));
    layer2_outputs(666) <= layer1_outputs(5128);
    layer2_outputs(667) <= not(layer1_outputs(4353));
    layer2_outputs(668) <= not((layer1_outputs(2124)) and (layer1_outputs(4781)));
    layer2_outputs(669) <= not(layer1_outputs(5215));
    layer2_outputs(670) <= layer1_outputs(2196);
    layer2_outputs(671) <= layer1_outputs(1898);
    layer2_outputs(672) <= '0';
    layer2_outputs(673) <= '0';
    layer2_outputs(674) <= layer1_outputs(7487);
    layer2_outputs(675) <= (layer1_outputs(2630)) and not (layer1_outputs(9836));
    layer2_outputs(676) <= (layer1_outputs(1987)) and not (layer1_outputs(3194));
    layer2_outputs(677) <= layer1_outputs(726);
    layer2_outputs(678) <= not(layer1_outputs(4307)) or (layer1_outputs(1701));
    layer2_outputs(679) <= layer1_outputs(2424);
    layer2_outputs(680) <= layer1_outputs(9185);
    layer2_outputs(681) <= layer1_outputs(201);
    layer2_outputs(682) <= layer1_outputs(3278);
    layer2_outputs(683) <= layer1_outputs(1531);
    layer2_outputs(684) <= layer1_outputs(8658);
    layer2_outputs(685) <= (layer1_outputs(3104)) xor (layer1_outputs(3505));
    layer2_outputs(686) <= not((layer1_outputs(10169)) or (layer1_outputs(5811)));
    layer2_outputs(687) <= (layer1_outputs(6511)) or (layer1_outputs(8151));
    layer2_outputs(688) <= layer1_outputs(671);
    layer2_outputs(689) <= not(layer1_outputs(9758));
    layer2_outputs(690) <= (layer1_outputs(7062)) and (layer1_outputs(9724));
    layer2_outputs(691) <= not(layer1_outputs(7719));
    layer2_outputs(692) <= not((layer1_outputs(4350)) or (layer1_outputs(6369)));
    layer2_outputs(693) <= not(layer1_outputs(215));
    layer2_outputs(694) <= layer1_outputs(1136);
    layer2_outputs(695) <= (layer1_outputs(4918)) and not (layer1_outputs(9319));
    layer2_outputs(696) <= layer1_outputs(4761);
    layer2_outputs(697) <= layer1_outputs(4700);
    layer2_outputs(698) <= not(layer1_outputs(9454)) or (layer1_outputs(2691));
    layer2_outputs(699) <= not(layer1_outputs(8170)) or (layer1_outputs(4905));
    layer2_outputs(700) <= layer1_outputs(679);
    layer2_outputs(701) <= '0';
    layer2_outputs(702) <= not((layer1_outputs(6839)) or (layer1_outputs(2169)));
    layer2_outputs(703) <= not(layer1_outputs(3628)) or (layer1_outputs(2423));
    layer2_outputs(704) <= not(layer1_outputs(2588));
    layer2_outputs(705) <= not(layer1_outputs(6753));
    layer2_outputs(706) <= (layer1_outputs(3898)) or (layer1_outputs(3896));
    layer2_outputs(707) <= not(layer1_outputs(6907));
    layer2_outputs(708) <= not(layer1_outputs(7990));
    layer2_outputs(709) <= layer1_outputs(6861);
    layer2_outputs(710) <= (layer1_outputs(5490)) and not (layer1_outputs(2467));
    layer2_outputs(711) <= (layer1_outputs(9140)) and not (layer1_outputs(7513));
    layer2_outputs(712) <= layer1_outputs(4514);
    layer2_outputs(713) <= layer1_outputs(5009);
    layer2_outputs(714) <= not(layer1_outputs(1747)) or (layer1_outputs(983));
    layer2_outputs(715) <= (layer1_outputs(4652)) and (layer1_outputs(3071));
    layer2_outputs(716) <= layer1_outputs(371);
    layer2_outputs(717) <= layer1_outputs(9552);
    layer2_outputs(718) <= not(layer1_outputs(5600));
    layer2_outputs(719) <= not((layer1_outputs(3544)) or (layer1_outputs(3207)));
    layer2_outputs(720) <= (layer1_outputs(5714)) and not (layer1_outputs(4325));
    layer2_outputs(721) <= layer1_outputs(5851);
    layer2_outputs(722) <= (layer1_outputs(8098)) or (layer1_outputs(1181));
    layer2_outputs(723) <= (layer1_outputs(3977)) and not (layer1_outputs(3253));
    layer2_outputs(724) <= not(layer1_outputs(3429));
    layer2_outputs(725) <= (layer1_outputs(5706)) or (layer1_outputs(6418));
    layer2_outputs(726) <= not((layer1_outputs(5147)) xor (layer1_outputs(7853)));
    layer2_outputs(727) <= '1';
    layer2_outputs(728) <= not(layer1_outputs(7780));
    layer2_outputs(729) <= (layer1_outputs(1191)) or (layer1_outputs(4297));
    layer2_outputs(730) <= not((layer1_outputs(4901)) or (layer1_outputs(2522)));
    layer2_outputs(731) <= (layer1_outputs(4715)) and (layer1_outputs(10207));
    layer2_outputs(732) <= not((layer1_outputs(2604)) or (layer1_outputs(4275)));
    layer2_outputs(733) <= not(layer1_outputs(6460)) or (layer1_outputs(4699));
    layer2_outputs(734) <= not((layer1_outputs(10185)) or (layer1_outputs(10115)));
    layer2_outputs(735) <= (layer1_outputs(2898)) or (layer1_outputs(5491));
    layer2_outputs(736) <= not(layer1_outputs(12));
    layer2_outputs(737) <= (layer1_outputs(1645)) xor (layer1_outputs(2695));
    layer2_outputs(738) <= layer1_outputs(4901);
    layer2_outputs(739) <= not((layer1_outputs(6222)) or (layer1_outputs(3269)));
    layer2_outputs(740) <= not((layer1_outputs(7561)) and (layer1_outputs(8933)));
    layer2_outputs(741) <= not(layer1_outputs(2981));
    layer2_outputs(742) <= (layer1_outputs(4024)) and not (layer1_outputs(9355));
    layer2_outputs(743) <= layer1_outputs(1936);
    layer2_outputs(744) <= '1';
    layer2_outputs(745) <= layer1_outputs(5038);
    layer2_outputs(746) <= layer1_outputs(4985);
    layer2_outputs(747) <= layer1_outputs(9815);
    layer2_outputs(748) <= layer1_outputs(3737);
    layer2_outputs(749) <= layer1_outputs(1720);
    layer2_outputs(750) <= (layer1_outputs(1753)) and (layer1_outputs(2226));
    layer2_outputs(751) <= '0';
    layer2_outputs(752) <= not((layer1_outputs(4850)) xor (layer1_outputs(241)));
    layer2_outputs(753) <= (layer1_outputs(9302)) and (layer1_outputs(5224));
    layer2_outputs(754) <= (layer1_outputs(7136)) and not (layer1_outputs(4982));
    layer2_outputs(755) <= layer1_outputs(4641);
    layer2_outputs(756) <= '1';
    layer2_outputs(757) <= (layer1_outputs(4508)) and not (layer1_outputs(2266));
    layer2_outputs(758) <= (layer1_outputs(4622)) and (layer1_outputs(1856));
    layer2_outputs(759) <= not(layer1_outputs(7859));
    layer2_outputs(760) <= layer1_outputs(10224);
    layer2_outputs(761) <= (layer1_outputs(2544)) and not (layer1_outputs(5069));
    layer2_outputs(762) <= (layer1_outputs(399)) or (layer1_outputs(8934));
    layer2_outputs(763) <= not((layer1_outputs(706)) and (layer1_outputs(4255)));
    layer2_outputs(764) <= (layer1_outputs(8357)) and not (layer1_outputs(560));
    layer2_outputs(765) <= not((layer1_outputs(4839)) xor (layer1_outputs(894)));
    layer2_outputs(766) <= not((layer1_outputs(10078)) or (layer1_outputs(9693)));
    layer2_outputs(767) <= layer1_outputs(55);
    layer2_outputs(768) <= (layer1_outputs(1016)) xor (layer1_outputs(8169));
    layer2_outputs(769) <= not((layer1_outputs(10128)) xor (layer1_outputs(4581)));
    layer2_outputs(770) <= not(layer1_outputs(2260));
    layer2_outputs(771) <= not(layer1_outputs(854)) or (layer1_outputs(10093));
    layer2_outputs(772) <= not(layer1_outputs(4865));
    layer2_outputs(773) <= layer1_outputs(9273);
    layer2_outputs(774) <= layer1_outputs(7208);
    layer2_outputs(775) <= (layer1_outputs(3476)) and not (layer1_outputs(7478));
    layer2_outputs(776) <= not((layer1_outputs(8697)) or (layer1_outputs(1686)));
    layer2_outputs(777) <= not(layer1_outputs(2628)) or (layer1_outputs(505));
    layer2_outputs(778) <= not(layer1_outputs(8524)) or (layer1_outputs(6209));
    layer2_outputs(779) <= not(layer1_outputs(1390));
    layer2_outputs(780) <= layer1_outputs(6050);
    layer2_outputs(781) <= not(layer1_outputs(187));
    layer2_outputs(782) <= not(layer1_outputs(7010));
    layer2_outputs(783) <= not(layer1_outputs(5631)) or (layer1_outputs(8611));
    layer2_outputs(784) <= not((layer1_outputs(7070)) xor (layer1_outputs(3894)));
    layer2_outputs(785) <= not((layer1_outputs(2555)) or (layer1_outputs(6132)));
    layer2_outputs(786) <= not(layer1_outputs(778));
    layer2_outputs(787) <= not(layer1_outputs(7856));
    layer2_outputs(788) <= layer1_outputs(6696);
    layer2_outputs(789) <= not((layer1_outputs(3538)) xor (layer1_outputs(4961)));
    layer2_outputs(790) <= layer1_outputs(408);
    layer2_outputs(791) <= (layer1_outputs(6710)) and not (layer1_outputs(5602));
    layer2_outputs(792) <= layer1_outputs(3267);
    layer2_outputs(793) <= layer1_outputs(589);
    layer2_outputs(794) <= not(layer1_outputs(9170));
    layer2_outputs(795) <= (layer1_outputs(2069)) and not (layer1_outputs(3569));
    layer2_outputs(796) <= layer1_outputs(183);
    layer2_outputs(797) <= (layer1_outputs(964)) or (layer1_outputs(5121));
    layer2_outputs(798) <= layer1_outputs(5106);
    layer2_outputs(799) <= not(layer1_outputs(8398)) or (layer1_outputs(7752));
    layer2_outputs(800) <= (layer1_outputs(3088)) or (layer1_outputs(3250));
    layer2_outputs(801) <= layer1_outputs(8409);
    layer2_outputs(802) <= not((layer1_outputs(6114)) and (layer1_outputs(3182)));
    layer2_outputs(803) <= (layer1_outputs(8046)) xor (layer1_outputs(2420));
    layer2_outputs(804) <= layer1_outputs(406);
    layer2_outputs(805) <= layer1_outputs(8542);
    layer2_outputs(806) <= layer1_outputs(5590);
    layer2_outputs(807) <= not(layer1_outputs(6883));
    layer2_outputs(808) <= (layer1_outputs(6983)) and not (layer1_outputs(1863));
    layer2_outputs(809) <= (layer1_outputs(8519)) and (layer1_outputs(7822));
    layer2_outputs(810) <= not(layer1_outputs(667));
    layer2_outputs(811) <= (layer1_outputs(8515)) or (layer1_outputs(2853));
    layer2_outputs(812) <= not(layer1_outputs(4025));
    layer2_outputs(813) <= layer1_outputs(4490);
    layer2_outputs(814) <= (layer1_outputs(5019)) and (layer1_outputs(7678));
    layer2_outputs(815) <= layer1_outputs(2546);
    layer2_outputs(816) <= not(layer1_outputs(3084)) or (layer1_outputs(3941));
    layer2_outputs(817) <= (layer1_outputs(8868)) xor (layer1_outputs(3148));
    layer2_outputs(818) <= (layer1_outputs(9017)) and (layer1_outputs(514));
    layer2_outputs(819) <= (layer1_outputs(5640)) or (layer1_outputs(6887));
    layer2_outputs(820) <= layer1_outputs(453);
    layer2_outputs(821) <= layer1_outputs(3708);
    layer2_outputs(822) <= not((layer1_outputs(2273)) and (layer1_outputs(21)));
    layer2_outputs(823) <= '1';
    layer2_outputs(824) <= not((layer1_outputs(3214)) or (layer1_outputs(1054)));
    layer2_outputs(825) <= not(layer1_outputs(4644));
    layer2_outputs(826) <= (layer1_outputs(1049)) and not (layer1_outputs(8225));
    layer2_outputs(827) <= layer1_outputs(9650);
    layer2_outputs(828) <= layer1_outputs(4679);
    layer2_outputs(829) <= (layer1_outputs(2675)) and not (layer1_outputs(8001));
    layer2_outputs(830) <= not((layer1_outputs(1499)) xor (layer1_outputs(8499)));
    layer2_outputs(831) <= not(layer1_outputs(6448));
    layer2_outputs(832) <= not(layer1_outputs(1132)) or (layer1_outputs(5812));
    layer2_outputs(833) <= not((layer1_outputs(5073)) and (layer1_outputs(629)));
    layer2_outputs(834) <= (layer1_outputs(9327)) xor (layer1_outputs(4005));
    layer2_outputs(835) <= not(layer1_outputs(5097));
    layer2_outputs(836) <= not((layer1_outputs(1931)) xor (layer1_outputs(4764)));
    layer2_outputs(837) <= (layer1_outputs(4634)) and (layer1_outputs(6123));
    layer2_outputs(838) <= not((layer1_outputs(8303)) xor (layer1_outputs(2544)));
    layer2_outputs(839) <= not(layer1_outputs(2663)) or (layer1_outputs(1301));
    layer2_outputs(840) <= (layer1_outputs(155)) xor (layer1_outputs(6642));
    layer2_outputs(841) <= (layer1_outputs(6173)) or (layer1_outputs(6848));
    layer2_outputs(842) <= (layer1_outputs(9876)) and not (layer1_outputs(2852));
    layer2_outputs(843) <= not((layer1_outputs(3973)) xor (layer1_outputs(7237)));
    layer2_outputs(844) <= (layer1_outputs(8498)) and not (layer1_outputs(8818));
    layer2_outputs(845) <= not(layer1_outputs(3937));
    layer2_outputs(846) <= not((layer1_outputs(643)) xor (layer1_outputs(1163)));
    layer2_outputs(847) <= not((layer1_outputs(6843)) xor (layer1_outputs(6281)));
    layer2_outputs(848) <= not((layer1_outputs(1924)) or (layer1_outputs(9674)));
    layer2_outputs(849) <= layer1_outputs(5277);
    layer2_outputs(850) <= layer1_outputs(222);
    layer2_outputs(851) <= (layer1_outputs(5392)) or (layer1_outputs(7784));
    layer2_outputs(852) <= layer1_outputs(7919);
    layer2_outputs(853) <= (layer1_outputs(6469)) xor (layer1_outputs(3107));
    layer2_outputs(854) <= not((layer1_outputs(1967)) or (layer1_outputs(2824)));
    layer2_outputs(855) <= layer1_outputs(4404);
    layer2_outputs(856) <= not(layer1_outputs(2186));
    layer2_outputs(857) <= layer1_outputs(6743);
    layer2_outputs(858) <= not(layer1_outputs(9720)) or (layer1_outputs(9456));
    layer2_outputs(859) <= not((layer1_outputs(7697)) and (layer1_outputs(5163)));
    layer2_outputs(860) <= (layer1_outputs(54)) xor (layer1_outputs(9528));
    layer2_outputs(861) <= layer1_outputs(5246);
    layer2_outputs(862) <= not(layer1_outputs(186));
    layer2_outputs(863) <= (layer1_outputs(892)) or (layer1_outputs(3771));
    layer2_outputs(864) <= layer1_outputs(1560);
    layer2_outputs(865) <= not((layer1_outputs(6921)) xor (layer1_outputs(3077)));
    layer2_outputs(866) <= not(layer1_outputs(1554));
    layer2_outputs(867) <= (layer1_outputs(5688)) and (layer1_outputs(9080));
    layer2_outputs(868) <= not(layer1_outputs(8695)) or (layer1_outputs(9941));
    layer2_outputs(869) <= not((layer1_outputs(3918)) xor (layer1_outputs(240)));
    layer2_outputs(870) <= layer1_outputs(1195);
    layer2_outputs(871) <= layer1_outputs(940);
    layer2_outputs(872) <= (layer1_outputs(6594)) xor (layer1_outputs(3521));
    layer2_outputs(873) <= (layer1_outputs(5169)) and not (layer1_outputs(1072));
    layer2_outputs(874) <= not((layer1_outputs(5808)) xor (layer1_outputs(7107)));
    layer2_outputs(875) <= not(layer1_outputs(8320)) or (layer1_outputs(2728));
    layer2_outputs(876) <= layer1_outputs(8148);
    layer2_outputs(877) <= (layer1_outputs(2719)) and not (layer1_outputs(7539));
    layer2_outputs(878) <= layer1_outputs(6231);
    layer2_outputs(879) <= not(layer1_outputs(9911));
    layer2_outputs(880) <= not(layer1_outputs(9317));
    layer2_outputs(881) <= not((layer1_outputs(7339)) and (layer1_outputs(8567)));
    layer2_outputs(882) <= not(layer1_outputs(8651));
    layer2_outputs(883) <= not(layer1_outputs(8506));
    layer2_outputs(884) <= not(layer1_outputs(7117));
    layer2_outputs(885) <= not((layer1_outputs(4896)) or (layer1_outputs(7188)));
    layer2_outputs(886) <= (layer1_outputs(4932)) and (layer1_outputs(3658));
    layer2_outputs(887) <= not(layer1_outputs(4115));
    layer2_outputs(888) <= not(layer1_outputs(2389));
    layer2_outputs(889) <= (layer1_outputs(2280)) xor (layer1_outputs(6292));
    layer2_outputs(890) <= not(layer1_outputs(6023)) or (layer1_outputs(5842));
    layer2_outputs(891) <= not(layer1_outputs(4919));
    layer2_outputs(892) <= layer1_outputs(4584);
    layer2_outputs(893) <= (layer1_outputs(10088)) xor (layer1_outputs(950));
    layer2_outputs(894) <= not(layer1_outputs(6044));
    layer2_outputs(895) <= not((layer1_outputs(1051)) and (layer1_outputs(5902)));
    layer2_outputs(896) <= not(layer1_outputs(2895)) or (layer1_outputs(5661));
    layer2_outputs(897) <= layer1_outputs(9554);
    layer2_outputs(898) <= not((layer1_outputs(5331)) and (layer1_outputs(6016)));
    layer2_outputs(899) <= layer1_outputs(8975);
    layer2_outputs(900) <= layer1_outputs(8020);
    layer2_outputs(901) <= not((layer1_outputs(114)) xor (layer1_outputs(5740)));
    layer2_outputs(902) <= not(layer1_outputs(3752));
    layer2_outputs(903) <= not(layer1_outputs(260));
    layer2_outputs(904) <= layer1_outputs(1805);
    layer2_outputs(905) <= (layer1_outputs(2040)) xor (layer1_outputs(8806));
    layer2_outputs(906) <= not(layer1_outputs(165));
    layer2_outputs(907) <= (layer1_outputs(8210)) xor (layer1_outputs(2398));
    layer2_outputs(908) <= not((layer1_outputs(8601)) xor (layer1_outputs(4940)));
    layer2_outputs(909) <= (layer1_outputs(353)) and not (layer1_outputs(9559));
    layer2_outputs(910) <= layer1_outputs(8434);
    layer2_outputs(911) <= not((layer1_outputs(3525)) or (layer1_outputs(2942)));
    layer2_outputs(912) <= layer1_outputs(1262);
    layer2_outputs(913) <= not(layer1_outputs(4166));
    layer2_outputs(914) <= (layer1_outputs(172)) xor (layer1_outputs(2418));
    layer2_outputs(915) <= not(layer1_outputs(7603)) or (layer1_outputs(2548));
    layer2_outputs(916) <= not(layer1_outputs(1844)) or (layer1_outputs(7371));
    layer2_outputs(917) <= not(layer1_outputs(8945)) or (layer1_outputs(9107));
    layer2_outputs(918) <= not((layer1_outputs(707)) and (layer1_outputs(4965)));
    layer2_outputs(919) <= layer1_outputs(4303);
    layer2_outputs(920) <= (layer1_outputs(3961)) and not (layer1_outputs(4394));
    layer2_outputs(921) <= not(layer1_outputs(4779)) or (layer1_outputs(2716));
    layer2_outputs(922) <= layer1_outputs(2960);
    layer2_outputs(923) <= (layer1_outputs(9006)) and (layer1_outputs(9723));
    layer2_outputs(924) <= layer1_outputs(6430);
    layer2_outputs(925) <= not((layer1_outputs(4663)) and (layer1_outputs(9088)));
    layer2_outputs(926) <= layer1_outputs(3602);
    layer2_outputs(927) <= (layer1_outputs(6103)) or (layer1_outputs(8001));
    layer2_outputs(928) <= not(layer1_outputs(5756));
    layer2_outputs(929) <= (layer1_outputs(1418)) and not (layer1_outputs(3153));
    layer2_outputs(930) <= not(layer1_outputs(5937));
    layer2_outputs(931) <= not(layer1_outputs(4911));
    layer2_outputs(932) <= not((layer1_outputs(4071)) xor (layer1_outputs(9804)));
    layer2_outputs(933) <= layer1_outputs(9871);
    layer2_outputs(934) <= layer1_outputs(7229);
    layer2_outputs(935) <= not((layer1_outputs(5680)) xor (layer1_outputs(2662)));
    layer2_outputs(936) <= not(layer1_outputs(2398)) or (layer1_outputs(6251));
    layer2_outputs(937) <= layer1_outputs(5593);
    layer2_outputs(938) <= not(layer1_outputs(7774));
    layer2_outputs(939) <= not(layer1_outputs(5402)) or (layer1_outputs(8919));
    layer2_outputs(940) <= not(layer1_outputs(5788));
    layer2_outputs(941) <= (layer1_outputs(10096)) and (layer1_outputs(2128));
    layer2_outputs(942) <= not((layer1_outputs(458)) and (layer1_outputs(3223)));
    layer2_outputs(943) <= (layer1_outputs(2290)) or (layer1_outputs(9063));
    layer2_outputs(944) <= not(layer1_outputs(8373));
    layer2_outputs(945) <= not(layer1_outputs(4140)) or (layer1_outputs(2710));
    layer2_outputs(946) <= layer1_outputs(7409);
    layer2_outputs(947) <= not(layer1_outputs(7981)) or (layer1_outputs(5077));
    layer2_outputs(948) <= '1';
    layer2_outputs(949) <= not(layer1_outputs(5999));
    layer2_outputs(950) <= not(layer1_outputs(56)) or (layer1_outputs(3038));
    layer2_outputs(951) <= '0';
    layer2_outputs(952) <= layer1_outputs(9840);
    layer2_outputs(953) <= not(layer1_outputs(2247));
    layer2_outputs(954) <= not((layer1_outputs(9198)) xor (layer1_outputs(5356)));
    layer2_outputs(955) <= not(layer1_outputs(5468));
    layer2_outputs(956) <= layer1_outputs(383);
    layer2_outputs(957) <= (layer1_outputs(7073)) or (layer1_outputs(1306));
    layer2_outputs(958) <= '1';
    layer2_outputs(959) <= layer1_outputs(6599);
    layer2_outputs(960) <= (layer1_outputs(737)) and not (layer1_outputs(295));
    layer2_outputs(961) <= (layer1_outputs(9020)) and not (layer1_outputs(6876));
    layer2_outputs(962) <= not((layer1_outputs(8368)) and (layer1_outputs(8697)));
    layer2_outputs(963) <= not((layer1_outputs(8494)) xor (layer1_outputs(3998)));
    layer2_outputs(964) <= not(layer1_outputs(7031)) or (layer1_outputs(1388));
    layer2_outputs(965) <= layer1_outputs(1609);
    layer2_outputs(966) <= layer1_outputs(8759);
    layer2_outputs(967) <= not((layer1_outputs(9571)) or (layer1_outputs(7806)));
    layer2_outputs(968) <= layer1_outputs(1885);
    layer2_outputs(969) <= not(layer1_outputs(8782));
    layer2_outputs(970) <= (layer1_outputs(8206)) and not (layer1_outputs(7313));
    layer2_outputs(971) <= (layer1_outputs(3236)) and not (layer1_outputs(8789));
    layer2_outputs(972) <= not(layer1_outputs(7345));
    layer2_outputs(973) <= not((layer1_outputs(6699)) xor (layer1_outputs(8072)));
    layer2_outputs(974) <= layer1_outputs(797);
    layer2_outputs(975) <= layer1_outputs(581);
    layer2_outputs(976) <= (layer1_outputs(8013)) or (layer1_outputs(336));
    layer2_outputs(977) <= not(layer1_outputs(9690));
    layer2_outputs(978) <= (layer1_outputs(1451)) or (layer1_outputs(5233));
    layer2_outputs(979) <= not((layer1_outputs(7291)) or (layer1_outputs(4556)));
    layer2_outputs(980) <= layer1_outputs(1697);
    layer2_outputs(981) <= layer1_outputs(120);
    layer2_outputs(982) <= (layer1_outputs(8477)) and not (layer1_outputs(2929));
    layer2_outputs(983) <= not(layer1_outputs(9029));
    layer2_outputs(984) <= not(layer1_outputs(5592));
    layer2_outputs(985) <= not((layer1_outputs(7963)) xor (layer1_outputs(7989)));
    layer2_outputs(986) <= (layer1_outputs(8095)) and not (layer1_outputs(2728));
    layer2_outputs(987) <= (layer1_outputs(9616)) and (layer1_outputs(1951));
    layer2_outputs(988) <= not((layer1_outputs(6976)) or (layer1_outputs(7772)));
    layer2_outputs(989) <= layer1_outputs(7443);
    layer2_outputs(990) <= (layer1_outputs(9201)) xor (layer1_outputs(7805));
    layer2_outputs(991) <= (layer1_outputs(8692)) and not (layer1_outputs(3630));
    layer2_outputs(992) <= (layer1_outputs(2402)) or (layer1_outputs(149));
    layer2_outputs(993) <= not(layer1_outputs(10010));
    layer2_outputs(994) <= (layer1_outputs(1273)) or (layer1_outputs(4295));
    layer2_outputs(995) <= layer1_outputs(7938);
    layer2_outputs(996) <= layer1_outputs(1341);
    layer2_outputs(997) <= layer1_outputs(6959);
    layer2_outputs(998) <= not((layer1_outputs(4324)) xor (layer1_outputs(6187)));
    layer2_outputs(999) <= not(layer1_outputs(9331)) or (layer1_outputs(6201));
    layer2_outputs(1000) <= layer1_outputs(6038);
    layer2_outputs(1001) <= layer1_outputs(5074);
    layer2_outputs(1002) <= not(layer1_outputs(5753));
    layer2_outputs(1003) <= layer1_outputs(8940);
    layer2_outputs(1004) <= layer1_outputs(4173);
    layer2_outputs(1005) <= not(layer1_outputs(1917));
    layer2_outputs(1006) <= layer1_outputs(5384);
    layer2_outputs(1007) <= not(layer1_outputs(1383)) or (layer1_outputs(8028));
    layer2_outputs(1008) <= not(layer1_outputs(8932));
    layer2_outputs(1009) <= (layer1_outputs(3106)) and not (layer1_outputs(1703));
    layer2_outputs(1010) <= not((layer1_outputs(8204)) xor (layer1_outputs(5511)));
    layer2_outputs(1011) <= (layer1_outputs(5542)) and not (layer1_outputs(7166));
    layer2_outputs(1012) <= layer1_outputs(4253);
    layer2_outputs(1013) <= (layer1_outputs(3410)) xor (layer1_outputs(1880));
    layer2_outputs(1014) <= (layer1_outputs(895)) and not (layer1_outputs(6685));
    layer2_outputs(1015) <= (layer1_outputs(7828)) or (layer1_outputs(6499));
    layer2_outputs(1016) <= '1';
    layer2_outputs(1017) <= (layer1_outputs(8225)) and not (layer1_outputs(770));
    layer2_outputs(1018) <= (layer1_outputs(10203)) xor (layer1_outputs(8536));
    layer2_outputs(1019) <= not(layer1_outputs(2709)) or (layer1_outputs(5223));
    layer2_outputs(1020) <= not(layer1_outputs(3004)) or (layer1_outputs(4537));
    layer2_outputs(1021) <= not(layer1_outputs(3504));
    layer2_outputs(1022) <= not(layer1_outputs(9763));
    layer2_outputs(1023) <= (layer1_outputs(1227)) and (layer1_outputs(9897));
    layer2_outputs(1024) <= (layer1_outputs(1721)) and not (layer1_outputs(4481));
    layer2_outputs(1025) <= layer1_outputs(5871);
    layer2_outputs(1026) <= not(layer1_outputs(2863));
    layer2_outputs(1027) <= not(layer1_outputs(6652));
    layer2_outputs(1028) <= not(layer1_outputs(2690)) or (layer1_outputs(2850));
    layer2_outputs(1029) <= not((layer1_outputs(1680)) or (layer1_outputs(2952)));
    layer2_outputs(1030) <= layer1_outputs(3023);
    layer2_outputs(1031) <= layer1_outputs(4413);
    layer2_outputs(1032) <= not(layer1_outputs(8029)) or (layer1_outputs(9562));
    layer2_outputs(1033) <= layer1_outputs(7543);
    layer2_outputs(1034) <= (layer1_outputs(1697)) and not (layer1_outputs(4560));
    layer2_outputs(1035) <= not(layer1_outputs(1966)) or (layer1_outputs(5867));
    layer2_outputs(1036) <= not(layer1_outputs(860));
    layer2_outputs(1037) <= not(layer1_outputs(3160));
    layer2_outputs(1038) <= not(layer1_outputs(2423));
    layer2_outputs(1039) <= (layer1_outputs(525)) and (layer1_outputs(4877));
    layer2_outputs(1040) <= not(layer1_outputs(974));
    layer2_outputs(1041) <= not((layer1_outputs(3259)) or (layer1_outputs(3373)));
    layer2_outputs(1042) <= (layer1_outputs(7915)) and (layer1_outputs(8825));
    layer2_outputs(1043) <= not((layer1_outputs(9737)) and (layer1_outputs(8474)));
    layer2_outputs(1044) <= not(layer1_outputs(9654));
    layer2_outputs(1045) <= layer1_outputs(9190);
    layer2_outputs(1046) <= layer1_outputs(2600);
    layer2_outputs(1047) <= not(layer1_outputs(365));
    layer2_outputs(1048) <= layer1_outputs(4623);
    layer2_outputs(1049) <= not((layer1_outputs(300)) and (layer1_outputs(9318)));
    layer2_outputs(1050) <= not(layer1_outputs(610));
    layer2_outputs(1051) <= not((layer1_outputs(3313)) xor (layer1_outputs(8634)));
    layer2_outputs(1052) <= not(layer1_outputs(1980)) or (layer1_outputs(6525));
    layer2_outputs(1053) <= (layer1_outputs(5435)) xor (layer1_outputs(6285));
    layer2_outputs(1054) <= layer1_outputs(9474);
    layer2_outputs(1055) <= not(layer1_outputs(4677)) or (layer1_outputs(3384));
    layer2_outputs(1056) <= not(layer1_outputs(2070));
    layer2_outputs(1057) <= not(layer1_outputs(8152));
    layer2_outputs(1058) <= (layer1_outputs(4355)) or (layer1_outputs(5912));
    layer2_outputs(1059) <= layer1_outputs(7814);
    layer2_outputs(1060) <= (layer1_outputs(9339)) xor (layer1_outputs(6110));
    layer2_outputs(1061) <= layer1_outputs(2405);
    layer2_outputs(1062) <= (layer1_outputs(5066)) and (layer1_outputs(4106));
    layer2_outputs(1063) <= not(layer1_outputs(1201));
    layer2_outputs(1064) <= layer1_outputs(2012);
    layer2_outputs(1065) <= not(layer1_outputs(7471));
    layer2_outputs(1066) <= not((layer1_outputs(2849)) or (layer1_outputs(374)));
    layer2_outputs(1067) <= '1';
    layer2_outputs(1068) <= not((layer1_outputs(6611)) xor (layer1_outputs(6810)));
    layer2_outputs(1069) <= not((layer1_outputs(4897)) and (layer1_outputs(3309)));
    layer2_outputs(1070) <= (layer1_outputs(5763)) and (layer1_outputs(491));
    layer2_outputs(1071) <= (layer1_outputs(3702)) and (layer1_outputs(6282));
    layer2_outputs(1072) <= (layer1_outputs(5230)) and not (layer1_outputs(6066));
    layer2_outputs(1073) <= (layer1_outputs(2756)) and not (layer1_outputs(8527));
    layer2_outputs(1074) <= layer1_outputs(3409);
    layer2_outputs(1075) <= (layer1_outputs(993)) and not (layer1_outputs(5414));
    layer2_outputs(1076) <= layer1_outputs(4694);
    layer2_outputs(1077) <= not((layer1_outputs(4669)) xor (layer1_outputs(8326)));
    layer2_outputs(1078) <= (layer1_outputs(3664)) and not (layer1_outputs(3763));
    layer2_outputs(1079) <= not(layer1_outputs(4359));
    layer2_outputs(1080) <= (layer1_outputs(7834)) and not (layer1_outputs(5802));
    layer2_outputs(1081) <= not((layer1_outputs(6228)) and (layer1_outputs(7740)));
    layer2_outputs(1082) <= (layer1_outputs(8837)) and (layer1_outputs(2643));
    layer2_outputs(1083) <= not(layer1_outputs(3482)) or (layer1_outputs(9564));
    layer2_outputs(1084) <= not((layer1_outputs(3454)) and (layer1_outputs(4783)));
    layer2_outputs(1085) <= layer1_outputs(1578);
    layer2_outputs(1086) <= (layer1_outputs(5300)) xor (layer1_outputs(7662));
    layer2_outputs(1087) <= layer1_outputs(2689);
    layer2_outputs(1088) <= (layer1_outputs(5931)) and not (layer1_outputs(3026));
    layer2_outputs(1089) <= (layer1_outputs(2134)) and (layer1_outputs(596));
    layer2_outputs(1090) <= not(layer1_outputs(661));
    layer2_outputs(1091) <= not((layer1_outputs(8550)) and (layer1_outputs(2261)));
    layer2_outputs(1092) <= (layer1_outputs(3677)) xor (layer1_outputs(2540));
    layer2_outputs(1093) <= not(layer1_outputs(7090));
    layer2_outputs(1094) <= not(layer1_outputs(5449));
    layer2_outputs(1095) <= (layer1_outputs(3731)) or (layer1_outputs(1259));
    layer2_outputs(1096) <= not((layer1_outputs(2653)) xor (layer1_outputs(8949)));
    layer2_outputs(1097) <= (layer1_outputs(9230)) and not (layer1_outputs(4687));
    layer2_outputs(1098) <= not(layer1_outputs(9068));
    layer2_outputs(1099) <= (layer1_outputs(6279)) and not (layer1_outputs(3016));
    layer2_outputs(1100) <= not(layer1_outputs(7934));
    layer2_outputs(1101) <= not(layer1_outputs(1449));
    layer2_outputs(1102) <= (layer1_outputs(1148)) and not (layer1_outputs(3169));
    layer2_outputs(1103) <= layer1_outputs(2108);
    layer2_outputs(1104) <= not(layer1_outputs(3956));
    layer2_outputs(1105) <= (layer1_outputs(9282)) or (layer1_outputs(2543));
    layer2_outputs(1106) <= not((layer1_outputs(4230)) or (layer1_outputs(6632)));
    layer2_outputs(1107) <= (layer1_outputs(410)) and not (layer1_outputs(8482));
    layer2_outputs(1108) <= not(layer1_outputs(1587)) or (layer1_outputs(9212));
    layer2_outputs(1109) <= (layer1_outputs(8944)) or (layer1_outputs(7373));
    layer2_outputs(1110) <= not(layer1_outputs(4515)) or (layer1_outputs(9146));
    layer2_outputs(1111) <= not(layer1_outputs(10044)) or (layer1_outputs(8801));
    layer2_outputs(1112) <= '0';
    layer2_outputs(1113) <= not((layer1_outputs(5791)) xor (layer1_outputs(5585)));
    layer2_outputs(1114) <= (layer1_outputs(9909)) xor (layer1_outputs(5769));
    layer2_outputs(1115) <= (layer1_outputs(5240)) and not (layer1_outputs(4223));
    layer2_outputs(1116) <= layer1_outputs(4408);
    layer2_outputs(1117) <= not(layer1_outputs(8512)) or (layer1_outputs(6666));
    layer2_outputs(1118) <= not(layer1_outputs(7892));
    layer2_outputs(1119) <= not(layer1_outputs(1596));
    layer2_outputs(1120) <= layer1_outputs(7522);
    layer2_outputs(1121) <= not(layer1_outputs(6655));
    layer2_outputs(1122) <= not(layer1_outputs(7724));
    layer2_outputs(1123) <= not(layer1_outputs(1913));
    layer2_outputs(1124) <= (layer1_outputs(279)) and not (layer1_outputs(4293));
    layer2_outputs(1125) <= not(layer1_outputs(4484));
    layer2_outputs(1126) <= (layer1_outputs(6094)) xor (layer1_outputs(9602));
    layer2_outputs(1127) <= (layer1_outputs(3402)) and not (layer1_outputs(2084));
    layer2_outputs(1128) <= '1';
    layer2_outputs(1129) <= not((layer1_outputs(2100)) and (layer1_outputs(3753)));
    layer2_outputs(1130) <= not((layer1_outputs(6391)) or (layer1_outputs(9092)));
    layer2_outputs(1131) <= (layer1_outputs(2922)) and not (layer1_outputs(8904));
    layer2_outputs(1132) <= layer1_outputs(3530);
    layer2_outputs(1133) <= '1';
    layer2_outputs(1134) <= (layer1_outputs(7849)) or (layer1_outputs(3850));
    layer2_outputs(1135) <= (layer1_outputs(10179)) or (layer1_outputs(5400));
    layer2_outputs(1136) <= layer1_outputs(10074);
    layer2_outputs(1137) <= not((layer1_outputs(8925)) and (layer1_outputs(1129)));
    layer2_outputs(1138) <= layer1_outputs(9660);
    layer2_outputs(1139) <= not(layer1_outputs(700)) or (layer1_outputs(5744));
    layer2_outputs(1140) <= not(layer1_outputs(6886));
    layer2_outputs(1141) <= not(layer1_outputs(8306));
    layer2_outputs(1142) <= layer1_outputs(8080);
    layer2_outputs(1143) <= (layer1_outputs(3871)) and not (layer1_outputs(9710));
    layer2_outputs(1144) <= not(layer1_outputs(4006));
    layer2_outputs(1145) <= not(layer1_outputs(9344)) or (layer1_outputs(4575));
    layer2_outputs(1146) <= not(layer1_outputs(2071));
    layer2_outputs(1147) <= layer1_outputs(980);
    layer2_outputs(1148) <= not(layer1_outputs(8139));
    layer2_outputs(1149) <= not(layer1_outputs(9158));
    layer2_outputs(1150) <= '0';
    layer2_outputs(1151) <= (layer1_outputs(6376)) and not (layer1_outputs(6774));
    layer2_outputs(1152) <= '0';
    layer2_outputs(1153) <= not((layer1_outputs(1407)) and (layer1_outputs(2329)));
    layer2_outputs(1154) <= not(layer1_outputs(1387)) or (layer1_outputs(2452));
    layer2_outputs(1155) <= not((layer1_outputs(9352)) xor (layer1_outputs(380)));
    layer2_outputs(1156) <= (layer1_outputs(2092)) or (layer1_outputs(7915));
    layer2_outputs(1157) <= (layer1_outputs(7446)) and not (layer1_outputs(4367));
    layer2_outputs(1158) <= (layer1_outputs(3660)) and not (layer1_outputs(3712));
    layer2_outputs(1159) <= not((layer1_outputs(2530)) xor (layer1_outputs(9316)));
    layer2_outputs(1160) <= (layer1_outputs(3563)) or (layer1_outputs(6832));
    layer2_outputs(1161) <= not(layer1_outputs(9876)) or (layer1_outputs(9765));
    layer2_outputs(1162) <= (layer1_outputs(7314)) xor (layer1_outputs(5425));
    layer2_outputs(1163) <= (layer1_outputs(8557)) xor (layer1_outputs(3345));
    layer2_outputs(1164) <= (layer1_outputs(5526)) and (layer1_outputs(6564));
    layer2_outputs(1165) <= layer1_outputs(7432);
    layer2_outputs(1166) <= layer1_outputs(7476);
    layer2_outputs(1167) <= layer1_outputs(5247);
    layer2_outputs(1168) <= not(layer1_outputs(2048));
    layer2_outputs(1169) <= not((layer1_outputs(480)) or (layer1_outputs(9732)));
    layer2_outputs(1170) <= (layer1_outputs(4244)) and not (layer1_outputs(3900));
    layer2_outputs(1171) <= not(layer1_outputs(1446));
    layer2_outputs(1172) <= not(layer1_outputs(2975)) or (layer1_outputs(181));
    layer2_outputs(1173) <= not((layer1_outputs(754)) xor (layer1_outputs(5189)));
    layer2_outputs(1174) <= not((layer1_outputs(4881)) xor (layer1_outputs(2485)));
    layer2_outputs(1175) <= not(layer1_outputs(2018));
    layer2_outputs(1176) <= (layer1_outputs(6656)) xor (layer1_outputs(1777));
    layer2_outputs(1177) <= (layer1_outputs(2212)) and (layer1_outputs(3451));
    layer2_outputs(1178) <= layer1_outputs(8341);
    layer2_outputs(1179) <= not((layer1_outputs(2228)) or (layer1_outputs(3156)));
    layer2_outputs(1180) <= not(layer1_outputs(6751)) or (layer1_outputs(7328));
    layer2_outputs(1181) <= (layer1_outputs(1274)) xor (layer1_outputs(3025));
    layer2_outputs(1182) <= layer1_outputs(8745);
    layer2_outputs(1183) <= not((layer1_outputs(3292)) and (layer1_outputs(4712)));
    layer2_outputs(1184) <= (layer1_outputs(9195)) xor (layer1_outputs(4086));
    layer2_outputs(1185) <= (layer1_outputs(5213)) xor (layer1_outputs(8912));
    layer2_outputs(1186) <= not(layer1_outputs(8217));
    layer2_outputs(1187) <= not(layer1_outputs(5024));
    layer2_outputs(1188) <= not(layer1_outputs(5363));
    layer2_outputs(1189) <= (layer1_outputs(348)) and not (layer1_outputs(7294));
    layer2_outputs(1190) <= (layer1_outputs(9151)) and (layer1_outputs(437));
    layer2_outputs(1191) <= not((layer1_outputs(7177)) xor (layer1_outputs(3026)));
    layer2_outputs(1192) <= (layer1_outputs(7383)) or (layer1_outputs(885));
    layer2_outputs(1193) <= not(layer1_outputs(5134));
    layer2_outputs(1194) <= not(layer1_outputs(3450));
    layer2_outputs(1195) <= not(layer1_outputs(9899));
    layer2_outputs(1196) <= (layer1_outputs(8996)) and not (layer1_outputs(4823));
    layer2_outputs(1197) <= layer1_outputs(2352);
    layer2_outputs(1198) <= not((layer1_outputs(2116)) xor (layer1_outputs(5207)));
    layer2_outputs(1199) <= (layer1_outputs(7175)) and (layer1_outputs(8464));
    layer2_outputs(1200) <= not(layer1_outputs(2831));
    layer2_outputs(1201) <= (layer1_outputs(5254)) and not (layer1_outputs(239));
    layer2_outputs(1202) <= not(layer1_outputs(8559));
    layer2_outputs(1203) <= not(layer1_outputs(3280));
    layer2_outputs(1204) <= not((layer1_outputs(767)) xor (layer1_outputs(4042)));
    layer2_outputs(1205) <= layer1_outputs(2392);
    layer2_outputs(1206) <= layer1_outputs(9863);
    layer2_outputs(1207) <= (layer1_outputs(5304)) xor (layer1_outputs(5587));
    layer2_outputs(1208) <= (layer1_outputs(7593)) xor (layer1_outputs(3684));
    layer2_outputs(1209) <= (layer1_outputs(2511)) and not (layer1_outputs(8557));
    layer2_outputs(1210) <= not((layer1_outputs(1055)) and (layer1_outputs(1598)));
    layer2_outputs(1211) <= not(layer1_outputs(4202));
    layer2_outputs(1212) <= layer1_outputs(4798);
    layer2_outputs(1213) <= (layer1_outputs(9249)) or (layer1_outputs(6241));
    layer2_outputs(1214) <= (layer1_outputs(5192)) or (layer1_outputs(217));
    layer2_outputs(1215) <= not(layer1_outputs(3649)) or (layer1_outputs(235));
    layer2_outputs(1216) <= layer1_outputs(6342);
    layer2_outputs(1217) <= not(layer1_outputs(9005)) or (layer1_outputs(7129));
    layer2_outputs(1218) <= not(layer1_outputs(1236));
    layer2_outputs(1219) <= not(layer1_outputs(1813)) or (layer1_outputs(6927));
    layer2_outputs(1220) <= (layer1_outputs(7456)) or (layer1_outputs(6219));
    layer2_outputs(1221) <= not(layer1_outputs(2440)) or (layer1_outputs(332));
    layer2_outputs(1222) <= (layer1_outputs(6040)) or (layer1_outputs(7014));
    layer2_outputs(1223) <= layer1_outputs(9048);
    layer2_outputs(1224) <= layer1_outputs(18);
    layer2_outputs(1225) <= not((layer1_outputs(709)) and (layer1_outputs(3068)));
    layer2_outputs(1226) <= layer1_outputs(8974);
    layer2_outputs(1227) <= not(layer1_outputs(7240)) or (layer1_outputs(3812));
    layer2_outputs(1228) <= not(layer1_outputs(4433)) or (layer1_outputs(8048));
    layer2_outputs(1229) <= not((layer1_outputs(373)) and (layer1_outputs(4016)));
    layer2_outputs(1230) <= not((layer1_outputs(9533)) xor (layer1_outputs(6139)));
    layer2_outputs(1231) <= not((layer1_outputs(5326)) or (layer1_outputs(3537)));
    layer2_outputs(1232) <= (layer1_outputs(4332)) and not (layer1_outputs(9410));
    layer2_outputs(1233) <= not(layer1_outputs(7731));
    layer2_outputs(1234) <= not((layer1_outputs(3989)) or (layer1_outputs(1137)));
    layer2_outputs(1235) <= not(layer1_outputs(6059));
    layer2_outputs(1236) <= not(layer1_outputs(7735));
    layer2_outputs(1237) <= (layer1_outputs(2257)) xor (layer1_outputs(3641));
    layer2_outputs(1238) <= layer1_outputs(5316);
    layer2_outputs(1239) <= layer1_outputs(6876);
    layer2_outputs(1240) <= not(layer1_outputs(6341));
    layer2_outputs(1241) <= layer1_outputs(5835);
    layer2_outputs(1242) <= not(layer1_outputs(5293)) or (layer1_outputs(460));
    layer2_outputs(1243) <= not((layer1_outputs(3698)) or (layer1_outputs(3827)));
    layer2_outputs(1244) <= not(layer1_outputs(394));
    layer2_outputs(1245) <= (layer1_outputs(3366)) and not (layer1_outputs(2794));
    layer2_outputs(1246) <= (layer1_outputs(1535)) xor (layer1_outputs(2763));
    layer2_outputs(1247) <= not((layer1_outputs(5769)) and (layer1_outputs(914)));
    layer2_outputs(1248) <= not(layer1_outputs(7461));
    layer2_outputs(1249) <= not(layer1_outputs(5238));
    layer2_outputs(1250) <= layer1_outputs(5581);
    layer2_outputs(1251) <= not((layer1_outputs(7306)) xor (layer1_outputs(8621)));
    layer2_outputs(1252) <= not(layer1_outputs(5877)) or (layer1_outputs(3725));
    layer2_outputs(1253) <= not(layer1_outputs(7139));
    layer2_outputs(1254) <= not(layer1_outputs(9071));
    layer2_outputs(1255) <= layer1_outputs(2391);
    layer2_outputs(1256) <= layer1_outputs(3339);
    layer2_outputs(1257) <= not(layer1_outputs(3303));
    layer2_outputs(1258) <= layer1_outputs(8986);
    layer2_outputs(1259) <= layer1_outputs(4126);
    layer2_outputs(1260) <= (layer1_outputs(9411)) and not (layer1_outputs(1023));
    layer2_outputs(1261) <= layer1_outputs(2838);
    layer2_outputs(1262) <= not(layer1_outputs(8100));
    layer2_outputs(1263) <= (layer1_outputs(3502)) xor (layer1_outputs(8762));
    layer2_outputs(1264) <= not((layer1_outputs(9926)) xor (layer1_outputs(1167)));
    layer2_outputs(1265) <= not(layer1_outputs(5442)) or (layer1_outputs(9554));
    layer2_outputs(1266) <= not((layer1_outputs(9106)) xor (layer1_outputs(1058)));
    layer2_outputs(1267) <= (layer1_outputs(7543)) and (layer1_outputs(3059));
    layer2_outputs(1268) <= not(layer1_outputs(2262));
    layer2_outputs(1269) <= layer1_outputs(8574);
    layer2_outputs(1270) <= not(layer1_outputs(4112));
    layer2_outputs(1271) <= not(layer1_outputs(3322)) or (layer1_outputs(4604));
    layer2_outputs(1272) <= not(layer1_outputs(2434));
    layer2_outputs(1273) <= not(layer1_outputs(9364)) or (layer1_outputs(1068));
    layer2_outputs(1274) <= not(layer1_outputs(4295));
    layer2_outputs(1275) <= not(layer1_outputs(6662)) or (layer1_outputs(6687));
    layer2_outputs(1276) <= not(layer1_outputs(1974));
    layer2_outputs(1277) <= not((layer1_outputs(7966)) and (layer1_outputs(6395)));
    layer2_outputs(1278) <= not((layer1_outputs(5696)) xor (layer1_outputs(4618)));
    layer2_outputs(1279) <= layer1_outputs(3361);
    layer2_outputs(1280) <= not(layer1_outputs(8684));
    layer2_outputs(1281) <= layer1_outputs(2427);
    layer2_outputs(1282) <= not(layer1_outputs(703));
    layer2_outputs(1283) <= not((layer1_outputs(2662)) or (layer1_outputs(5795)));
    layer2_outputs(1284) <= layer1_outputs(5114);
    layer2_outputs(1285) <= not(layer1_outputs(8127));
    layer2_outputs(1286) <= (layer1_outputs(5779)) and (layer1_outputs(3560));
    layer2_outputs(1287) <= not((layer1_outputs(8658)) xor (layer1_outputs(1266)));
    layer2_outputs(1288) <= (layer1_outputs(3967)) xor (layer1_outputs(7535));
    layer2_outputs(1289) <= layer1_outputs(110);
    layer2_outputs(1290) <= layer1_outputs(5965);
    layer2_outputs(1291) <= (layer1_outputs(8799)) xor (layer1_outputs(9795));
    layer2_outputs(1292) <= (layer1_outputs(4277)) and not (layer1_outputs(2611));
    layer2_outputs(1293) <= (layer1_outputs(4962)) or (layer1_outputs(5148));
    layer2_outputs(1294) <= (layer1_outputs(1562)) and not (layer1_outputs(2784));
    layer2_outputs(1295) <= layer1_outputs(425);
    layer2_outputs(1296) <= layer1_outputs(1260);
    layer2_outputs(1297) <= (layer1_outputs(5429)) and (layer1_outputs(9167));
    layer2_outputs(1298) <= not(layer1_outputs(996));
    layer2_outputs(1299) <= not(layer1_outputs(4089));
    layer2_outputs(1300) <= not(layer1_outputs(5470)) or (layer1_outputs(9132));
    layer2_outputs(1301) <= not(layer1_outputs(4005));
    layer2_outputs(1302) <= (layer1_outputs(6776)) and not (layer1_outputs(1774));
    layer2_outputs(1303) <= (layer1_outputs(670)) or (layer1_outputs(728));
    layer2_outputs(1304) <= not(layer1_outputs(5582));
    layer2_outputs(1305) <= (layer1_outputs(8548)) xor (layer1_outputs(1116));
    layer2_outputs(1306) <= not(layer1_outputs(7645));
    layer2_outputs(1307) <= not(layer1_outputs(7017));
    layer2_outputs(1308) <= not((layer1_outputs(1606)) xor (layer1_outputs(7151)));
    layer2_outputs(1309) <= layer1_outputs(6120);
    layer2_outputs(1310) <= (layer1_outputs(3930)) xor (layer1_outputs(840));
    layer2_outputs(1311) <= (layer1_outputs(1797)) and not (layer1_outputs(915));
    layer2_outputs(1312) <= layer1_outputs(2432);
    layer2_outputs(1313) <= not((layer1_outputs(6466)) and (layer1_outputs(3811)));
    layer2_outputs(1314) <= layer1_outputs(4073);
    layer2_outputs(1315) <= layer1_outputs(2001);
    layer2_outputs(1316) <= layer1_outputs(9938);
    layer2_outputs(1317) <= not((layer1_outputs(9967)) xor (layer1_outputs(2656)));
    layer2_outputs(1318) <= layer1_outputs(7320);
    layer2_outputs(1319) <= not((layer1_outputs(8643)) or (layer1_outputs(2232)));
    layer2_outputs(1320) <= layer1_outputs(2906);
    layer2_outputs(1321) <= layer1_outputs(1300);
    layer2_outputs(1322) <= layer1_outputs(2148);
    layer2_outputs(1323) <= not(layer1_outputs(15));
    layer2_outputs(1324) <= (layer1_outputs(8633)) and (layer1_outputs(3100));
    layer2_outputs(1325) <= layer1_outputs(2548);
    layer2_outputs(1326) <= (layer1_outputs(1683)) and (layer1_outputs(2944));
    layer2_outputs(1327) <= not(layer1_outputs(6026)) or (layer1_outputs(3919));
    layer2_outputs(1328) <= layer1_outputs(6889);
    layer2_outputs(1329) <= layer1_outputs(8730);
    layer2_outputs(1330) <= (layer1_outputs(8260)) or (layer1_outputs(2322));
    layer2_outputs(1331) <= not(layer1_outputs(7582)) or (layer1_outputs(3908));
    layer2_outputs(1332) <= (layer1_outputs(1290)) or (layer1_outputs(3140));
    layer2_outputs(1333) <= (layer1_outputs(6506)) xor (layer1_outputs(2009));
    layer2_outputs(1334) <= (layer1_outputs(8706)) and not (layer1_outputs(705));
    layer2_outputs(1335) <= (layer1_outputs(3675)) or (layer1_outputs(4027));
    layer2_outputs(1336) <= layer1_outputs(4384);
    layer2_outputs(1337) <= not(layer1_outputs(2958));
    layer2_outputs(1338) <= not(layer1_outputs(4099));
    layer2_outputs(1339) <= (layer1_outputs(4864)) and (layer1_outputs(8404));
    layer2_outputs(1340) <= (layer1_outputs(6411)) and not (layer1_outputs(9735));
    layer2_outputs(1341) <= not(layer1_outputs(2811)) or (layer1_outputs(9803));
    layer2_outputs(1342) <= '0';
    layer2_outputs(1343) <= not((layer1_outputs(5596)) or (layer1_outputs(405)));
    layer2_outputs(1344) <= not(layer1_outputs(5246));
    layer2_outputs(1345) <= not((layer1_outputs(5533)) and (layer1_outputs(3197)));
    layer2_outputs(1346) <= not((layer1_outputs(4104)) and (layer1_outputs(1516)));
    layer2_outputs(1347) <= (layer1_outputs(9075)) or (layer1_outputs(2569));
    layer2_outputs(1348) <= (layer1_outputs(9860)) and not (layer1_outputs(9708));
    layer2_outputs(1349) <= not(layer1_outputs(9133));
    layer2_outputs(1350) <= not(layer1_outputs(6301));
    layer2_outputs(1351) <= (layer1_outputs(1144)) and not (layer1_outputs(6446));
    layer2_outputs(1352) <= layer1_outputs(9411);
    layer2_outputs(1353) <= not(layer1_outputs(520)) or (layer1_outputs(3905));
    layer2_outputs(1354) <= layer1_outputs(8047);
    layer2_outputs(1355) <= layer1_outputs(1818);
    layer2_outputs(1356) <= not(layer1_outputs(9245));
    layer2_outputs(1357) <= not(layer1_outputs(4497));
    layer2_outputs(1358) <= layer1_outputs(7763);
    layer2_outputs(1359) <= not(layer1_outputs(270));
    layer2_outputs(1360) <= (layer1_outputs(1930)) and not (layer1_outputs(6095));
    layer2_outputs(1361) <= layer1_outputs(6002);
    layer2_outputs(1362) <= not((layer1_outputs(8139)) xor (layer1_outputs(5471)));
    layer2_outputs(1363) <= not((layer1_outputs(9950)) or (layer1_outputs(2776)));
    layer2_outputs(1364) <= layer1_outputs(3137);
    layer2_outputs(1365) <= layer1_outputs(384);
    layer2_outputs(1366) <= not(layer1_outputs(741)) or (layer1_outputs(9220));
    layer2_outputs(1367) <= not((layer1_outputs(5870)) xor (layer1_outputs(9710)));
    layer2_outputs(1368) <= not(layer1_outputs(7187));
    layer2_outputs(1369) <= not((layer1_outputs(3164)) xor (layer1_outputs(9166)));
    layer2_outputs(1370) <= (layer1_outputs(5390)) and not (layer1_outputs(5747));
    layer2_outputs(1371) <= (layer1_outputs(4394)) or (layer1_outputs(6576));
    layer2_outputs(1372) <= not(layer1_outputs(1846)) or (layer1_outputs(175));
    layer2_outputs(1373) <= layer1_outputs(9245);
    layer2_outputs(1374) <= layer1_outputs(2487);
    layer2_outputs(1375) <= layer1_outputs(7809);
    layer2_outputs(1376) <= (layer1_outputs(7672)) xor (layer1_outputs(8898));
    layer2_outputs(1377) <= not(layer1_outputs(9896));
    layer2_outputs(1378) <= not(layer1_outputs(4063));
    layer2_outputs(1379) <= not((layer1_outputs(1643)) xor (layer1_outputs(9126)));
    layer2_outputs(1380) <= layer1_outputs(1450);
    layer2_outputs(1381) <= layer1_outputs(8850);
    layer2_outputs(1382) <= (layer1_outputs(2517)) and not (layer1_outputs(4624));
    layer2_outputs(1383) <= not((layer1_outputs(8782)) and (layer1_outputs(7462)));
    layer2_outputs(1384) <= not(layer1_outputs(10027)) or (layer1_outputs(4650));
    layer2_outputs(1385) <= layer1_outputs(617);
    layer2_outputs(1386) <= (layer1_outputs(8363)) and (layer1_outputs(7715));
    layer2_outputs(1387) <= (layer1_outputs(6702)) and (layer1_outputs(4628));
    layer2_outputs(1388) <= not(layer1_outputs(7069));
    layer2_outputs(1389) <= (layer1_outputs(2707)) xor (layer1_outputs(6235));
    layer2_outputs(1390) <= not(layer1_outputs(7316));
    layer2_outputs(1391) <= not(layer1_outputs(7301));
    layer2_outputs(1392) <= not((layer1_outputs(8158)) or (layer1_outputs(6734)));
    layer2_outputs(1393) <= not(layer1_outputs(8800)) or (layer1_outputs(979));
    layer2_outputs(1394) <= (layer1_outputs(3761)) xor (layer1_outputs(5741));
    layer2_outputs(1395) <= not(layer1_outputs(6659));
    layer2_outputs(1396) <= '1';
    layer2_outputs(1397) <= not(layer1_outputs(9495));
    layer2_outputs(1398) <= layer1_outputs(5604);
    layer2_outputs(1399) <= not(layer1_outputs(148)) or (layer1_outputs(6637));
    layer2_outputs(1400) <= layer1_outputs(9728);
    layer2_outputs(1401) <= not(layer1_outputs(1830));
    layer2_outputs(1402) <= layer1_outputs(1872);
    layer2_outputs(1403) <= not((layer1_outputs(3935)) and (layer1_outputs(6512)));
    layer2_outputs(1404) <= layer1_outputs(33);
    layer2_outputs(1405) <= layer1_outputs(1337);
    layer2_outputs(1406) <= not(layer1_outputs(204));
    layer2_outputs(1407) <= not((layer1_outputs(2522)) xor (layer1_outputs(1998)));
    layer2_outputs(1408) <= layer1_outputs(2809);
    layer2_outputs(1409) <= not((layer1_outputs(2974)) and (layer1_outputs(4216)));
    layer2_outputs(1410) <= not(layer1_outputs(9620));
    layer2_outputs(1411) <= not((layer1_outputs(10239)) and (layer1_outputs(292)));
    layer2_outputs(1412) <= not(layer1_outputs(2007)) or (layer1_outputs(8182));
    layer2_outputs(1413) <= layer1_outputs(2880);
    layer2_outputs(1414) <= not(layer1_outputs(6274));
    layer2_outputs(1415) <= layer1_outputs(9178);
    layer2_outputs(1416) <= (layer1_outputs(8248)) or (layer1_outputs(1579));
    layer2_outputs(1417) <= layer1_outputs(1704);
    layer2_outputs(1418) <= layer1_outputs(576);
    layer2_outputs(1419) <= (layer1_outputs(5090)) and (layer1_outputs(8800));
    layer2_outputs(1420) <= not(layer1_outputs(8950));
    layer2_outputs(1421) <= not(layer1_outputs(3833));
    layer2_outputs(1422) <= not(layer1_outputs(4795)) or (layer1_outputs(10206));
    layer2_outputs(1423) <= layer1_outputs(9106);
    layer2_outputs(1424) <= not(layer1_outputs(2825));
    layer2_outputs(1425) <= layer1_outputs(5433);
    layer2_outputs(1426) <= layer1_outputs(1709);
    layer2_outputs(1427) <= not((layer1_outputs(2915)) xor (layer1_outputs(8585)));
    layer2_outputs(1428) <= layer1_outputs(6923);
    layer2_outputs(1429) <= not(layer1_outputs(6233));
    layer2_outputs(1430) <= not(layer1_outputs(383));
    layer2_outputs(1431) <= not(layer1_outputs(8356));
    layer2_outputs(1432) <= layer1_outputs(9415);
    layer2_outputs(1433) <= (layer1_outputs(950)) and not (layer1_outputs(9295));
    layer2_outputs(1434) <= not(layer1_outputs(7574));
    layer2_outputs(1435) <= not((layer1_outputs(1126)) and (layer1_outputs(6155)));
    layer2_outputs(1436) <= not((layer1_outputs(9969)) and (layer1_outputs(1064)));
    layer2_outputs(1437) <= (layer1_outputs(10046)) and not (layer1_outputs(5937));
    layer2_outputs(1438) <= not(layer1_outputs(4120));
    layer2_outputs(1439) <= not(layer1_outputs(9203));
    layer2_outputs(1440) <= not((layer1_outputs(1630)) and (layer1_outputs(4195)));
    layer2_outputs(1441) <= not(layer1_outputs(2049));
    layer2_outputs(1442) <= (layer1_outputs(9634)) xor (layer1_outputs(1927));
    layer2_outputs(1443) <= not(layer1_outputs(5748));
    layer2_outputs(1444) <= not(layer1_outputs(9682)) or (layer1_outputs(2627));
    layer2_outputs(1445) <= not((layer1_outputs(8530)) or (layer1_outputs(974)));
    layer2_outputs(1446) <= (layer1_outputs(1798)) or (layer1_outputs(5368));
    layer2_outputs(1447) <= not(layer1_outputs(2815)) or (layer1_outputs(1097));
    layer2_outputs(1448) <= not(layer1_outputs(8323)) or (layer1_outputs(4116));
    layer2_outputs(1449) <= (layer1_outputs(310)) and not (layer1_outputs(2602));
    layer2_outputs(1450) <= (layer1_outputs(5409)) and not (layer1_outputs(1625));
    layer2_outputs(1451) <= not(layer1_outputs(7098)) or (layer1_outputs(9227));
    layer2_outputs(1452) <= layer1_outputs(8484);
    layer2_outputs(1453) <= (layer1_outputs(1816)) xor (layer1_outputs(4780));
    layer2_outputs(1454) <= not(layer1_outputs(6867));
    layer2_outputs(1455) <= (layer1_outputs(8835)) and not (layer1_outputs(4504));
    layer2_outputs(1456) <= not(layer1_outputs(389));
    layer2_outputs(1457) <= not(layer1_outputs(7946));
    layer2_outputs(1458) <= (layer1_outputs(1250)) and not (layer1_outputs(1288));
    layer2_outputs(1459) <= not((layer1_outputs(1060)) xor (layer1_outputs(9375)));
    layer2_outputs(1460) <= not(layer1_outputs(7164));
    layer2_outputs(1461) <= not(layer1_outputs(9610)) or (layer1_outputs(8717));
    layer2_outputs(1462) <= not(layer1_outputs(10074));
    layer2_outputs(1463) <= not(layer1_outputs(3221));
    layer2_outputs(1464) <= not((layer1_outputs(4994)) xor (layer1_outputs(1628)));
    layer2_outputs(1465) <= not((layer1_outputs(2292)) xor (layer1_outputs(4605)));
    layer2_outputs(1466) <= (layer1_outputs(3533)) xor (layer1_outputs(5782));
    layer2_outputs(1467) <= not(layer1_outputs(9651)) or (layer1_outputs(5981));
    layer2_outputs(1468) <= not(layer1_outputs(3362)) or (layer1_outputs(9338));
    layer2_outputs(1469) <= not(layer1_outputs(5911));
    layer2_outputs(1470) <= not(layer1_outputs(2919));
    layer2_outputs(1471) <= not(layer1_outputs(1606));
    layer2_outputs(1472) <= (layer1_outputs(2595)) and (layer1_outputs(2185));
    layer2_outputs(1473) <= not(layer1_outputs(3756));
    layer2_outputs(1474) <= (layer1_outputs(5338)) and not (layer1_outputs(6616));
    layer2_outputs(1475) <= not(layer1_outputs(4732)) or (layer1_outputs(6290));
    layer2_outputs(1476) <= not(layer1_outputs(5541));
    layer2_outputs(1477) <= not(layer1_outputs(9319));
    layer2_outputs(1478) <= not(layer1_outputs(2965));
    layer2_outputs(1479) <= not((layer1_outputs(7521)) xor (layer1_outputs(1672)));
    layer2_outputs(1480) <= layer1_outputs(3660);
    layer2_outputs(1481) <= not(layer1_outputs(6133));
    layer2_outputs(1482) <= not(layer1_outputs(1958)) or (layer1_outputs(7728));
    layer2_outputs(1483) <= not((layer1_outputs(5005)) xor (layer1_outputs(9265)));
    layer2_outputs(1484) <= layer1_outputs(4887);
    layer2_outputs(1485) <= layer1_outputs(1325);
    layer2_outputs(1486) <= not((layer1_outputs(2167)) or (layer1_outputs(9905)));
    layer2_outputs(1487) <= not((layer1_outputs(6578)) or (layer1_outputs(948)));
    layer2_outputs(1488) <= not(layer1_outputs(5222));
    layer2_outputs(1489) <= not(layer1_outputs(6459));
    layer2_outputs(1490) <= not(layer1_outputs(1346)) or (layer1_outputs(2121));
    layer2_outputs(1491) <= not(layer1_outputs(5442));
    layer2_outputs(1492) <= (layer1_outputs(6004)) xor (layer1_outputs(7948));
    layer2_outputs(1493) <= not(layer1_outputs(9682));
    layer2_outputs(1494) <= not((layer1_outputs(8872)) and (layer1_outputs(4511)));
    layer2_outputs(1495) <= '0';
    layer2_outputs(1496) <= (layer1_outputs(2364)) and not (layer1_outputs(5334));
    layer2_outputs(1497) <= not(layer1_outputs(2594)) or (layer1_outputs(9214));
    layer2_outputs(1498) <= layer1_outputs(467);
    layer2_outputs(1499) <= (layer1_outputs(3794)) or (layer1_outputs(6962));
    layer2_outputs(1500) <= layer1_outputs(8494);
    layer2_outputs(1501) <= (layer1_outputs(7303)) xor (layer1_outputs(370));
    layer2_outputs(1502) <= not(layer1_outputs(3470));
    layer2_outputs(1503) <= '1';
    layer2_outputs(1504) <= not(layer1_outputs(2480)) or (layer1_outputs(3776));
    layer2_outputs(1505) <= not(layer1_outputs(7347));
    layer2_outputs(1506) <= layer1_outputs(1682);
    layer2_outputs(1507) <= (layer1_outputs(3907)) xor (layer1_outputs(1848));
    layer2_outputs(1508) <= not(layer1_outputs(4000)) or (layer1_outputs(8267));
    layer2_outputs(1509) <= layer1_outputs(8592);
    layer2_outputs(1510) <= layer1_outputs(488);
    layer2_outputs(1511) <= not(layer1_outputs(1406));
    layer2_outputs(1512) <= not(layer1_outputs(5460));
    layer2_outputs(1513) <= not((layer1_outputs(8598)) xor (layer1_outputs(986)));
    layer2_outputs(1514) <= (layer1_outputs(9091)) and not (layer1_outputs(2034));
    layer2_outputs(1515) <= not((layer1_outputs(6793)) and (layer1_outputs(1347)));
    layer2_outputs(1516) <= not(layer1_outputs(118));
    layer2_outputs(1517) <= not((layer1_outputs(2333)) xor (layer1_outputs(6635)));
    layer2_outputs(1518) <= layer1_outputs(2053);
    layer2_outputs(1519) <= not((layer1_outputs(4319)) xor (layer1_outputs(8471)));
    layer2_outputs(1520) <= not(layer1_outputs(1088)) or (layer1_outputs(7477));
    layer2_outputs(1521) <= (layer1_outputs(6905)) and (layer1_outputs(2462));
    layer2_outputs(1522) <= not(layer1_outputs(8273)) or (layer1_outputs(7206));
    layer2_outputs(1523) <= not(layer1_outputs(4528));
    layer2_outputs(1524) <= (layer1_outputs(3692)) or (layer1_outputs(1476));
    layer2_outputs(1525) <= not(layer1_outputs(2580)) or (layer1_outputs(3290));
    layer2_outputs(1526) <= not((layer1_outputs(5481)) xor (layer1_outputs(792)));
    layer2_outputs(1527) <= not(layer1_outputs(8927));
    layer2_outputs(1528) <= not(layer1_outputs(4056));
    layer2_outputs(1529) <= not(layer1_outputs(9790));
    layer2_outputs(1530) <= layer1_outputs(7495);
    layer2_outputs(1531) <= not((layer1_outputs(1204)) xor (layer1_outputs(9535)));
    layer2_outputs(1532) <= not((layer1_outputs(9638)) xor (layer1_outputs(9308)));
    layer2_outputs(1533) <= not(layer1_outputs(1166));
    layer2_outputs(1534) <= (layer1_outputs(8619)) and (layer1_outputs(3631));
    layer2_outputs(1535) <= layer1_outputs(6246);
    layer2_outputs(1536) <= not(layer1_outputs(7465));
    layer2_outputs(1537) <= not(layer1_outputs(1855)) or (layer1_outputs(6455));
    layer2_outputs(1538) <= layer1_outputs(6502);
    layer2_outputs(1539) <= not(layer1_outputs(10034)) or (layer1_outputs(4908));
    layer2_outputs(1540) <= layer1_outputs(9882);
    layer2_outputs(1541) <= not((layer1_outputs(10001)) and (layer1_outputs(6349)));
    layer2_outputs(1542) <= (layer1_outputs(6552)) and not (layer1_outputs(2249));
    layer2_outputs(1543) <= not(layer1_outputs(8785)) or (layer1_outputs(5163));
    layer2_outputs(1544) <= layer1_outputs(4792);
    layer2_outputs(1545) <= layer1_outputs(6753);
    layer2_outputs(1546) <= not(layer1_outputs(4260));
    layer2_outputs(1547) <= not(layer1_outputs(9853)) or (layer1_outputs(130));
    layer2_outputs(1548) <= not(layer1_outputs(7433));
    layer2_outputs(1549) <= not((layer1_outputs(938)) and (layer1_outputs(6177)));
    layer2_outputs(1550) <= (layer1_outputs(6223)) and not (layer1_outputs(6520));
    layer2_outputs(1551) <= not(layer1_outputs(2633)) or (layer1_outputs(7688));
    layer2_outputs(1552) <= layer1_outputs(9404);
    layer2_outputs(1553) <= (layer1_outputs(1735)) and not (layer1_outputs(3263));
    layer2_outputs(1554) <= not((layer1_outputs(6478)) xor (layer1_outputs(3922)));
    layer2_outputs(1555) <= (layer1_outputs(8962)) and not (layer1_outputs(3844));
    layer2_outputs(1556) <= not(layer1_outputs(4411));
    layer2_outputs(1557) <= layer1_outputs(3703);
    layer2_outputs(1558) <= layer1_outputs(2178);
    layer2_outputs(1559) <= layer1_outputs(2672);
    layer2_outputs(1560) <= not(layer1_outputs(8071));
    layer2_outputs(1561) <= not(layer1_outputs(5755));
    layer2_outputs(1562) <= layer1_outputs(1310);
    layer2_outputs(1563) <= (layer1_outputs(384)) and not (layer1_outputs(2532));
    layer2_outputs(1564) <= (layer1_outputs(9262)) and not (layer1_outputs(10153));
    layer2_outputs(1565) <= not((layer1_outputs(742)) and (layer1_outputs(6613)));
    layer2_outputs(1566) <= layer1_outputs(6515);
    layer2_outputs(1567) <= (layer1_outputs(7456)) or (layer1_outputs(6534));
    layer2_outputs(1568) <= not(layer1_outputs(9107));
    layer2_outputs(1569) <= not(layer1_outputs(1810));
    layer2_outputs(1570) <= layer1_outputs(8687);
    layer2_outputs(1571) <= layer1_outputs(1919);
    layer2_outputs(1572) <= not((layer1_outputs(5862)) or (layer1_outputs(5709)));
    layer2_outputs(1573) <= layer1_outputs(3654);
    layer2_outputs(1574) <= (layer1_outputs(10077)) and (layer1_outputs(552));
    layer2_outputs(1575) <= not(layer1_outputs(9512)) or (layer1_outputs(4360));
    layer2_outputs(1576) <= not(layer1_outputs(5819));
    layer2_outputs(1577) <= not(layer1_outputs(10071)) or (layer1_outputs(3294));
    layer2_outputs(1578) <= not(layer1_outputs(8901));
    layer2_outputs(1579) <= (layer1_outputs(3103)) xor (layer1_outputs(3162));
    layer2_outputs(1580) <= not(layer1_outputs(7195));
    layer2_outputs(1581) <= layer1_outputs(704);
    layer2_outputs(1582) <= not(layer1_outputs(3399));
    layer2_outputs(1583) <= not(layer1_outputs(2817)) or (layer1_outputs(4736));
    layer2_outputs(1584) <= '1';
    layer2_outputs(1585) <= (layer1_outputs(2210)) or (layer1_outputs(849));
    layer2_outputs(1586) <= (layer1_outputs(5946)) xor (layer1_outputs(7484));
    layer2_outputs(1587) <= layer1_outputs(2066);
    layer2_outputs(1588) <= not(layer1_outputs(5581));
    layer2_outputs(1589) <= (layer1_outputs(1270)) and not (layer1_outputs(5517));
    layer2_outputs(1590) <= not(layer1_outputs(719)) or (layer1_outputs(780));
    layer2_outputs(1591) <= layer1_outputs(2669);
    layer2_outputs(1592) <= not(layer1_outputs(8938));
    layer2_outputs(1593) <= layer1_outputs(8309);
    layer2_outputs(1594) <= not((layer1_outputs(3392)) xor (layer1_outputs(3499)));
    layer2_outputs(1595) <= layer1_outputs(2671);
    layer2_outputs(1596) <= (layer1_outputs(2986)) or (layer1_outputs(9705));
    layer2_outputs(1597) <= layer1_outputs(6722);
    layer2_outputs(1598) <= (layer1_outputs(9064)) and not (layer1_outputs(8290));
    layer2_outputs(1599) <= not(layer1_outputs(947));
    layer2_outputs(1600) <= not(layer1_outputs(6048));
    layer2_outputs(1601) <= not(layer1_outputs(8703)) or (layer1_outputs(8975));
    layer2_outputs(1602) <= not((layer1_outputs(869)) and (layer1_outputs(3463)));
    layer2_outputs(1603) <= not(layer1_outputs(4946));
    layer2_outputs(1604) <= not((layer1_outputs(554)) or (layer1_outputs(1043)));
    layer2_outputs(1605) <= layer1_outputs(656);
    layer2_outputs(1606) <= (layer1_outputs(7126)) or (layer1_outputs(3480));
    layer2_outputs(1607) <= layer1_outputs(6524);
    layer2_outputs(1608) <= not(layer1_outputs(7022));
    layer2_outputs(1609) <= not(layer1_outputs(8056)) or (layer1_outputs(7477));
    layer2_outputs(1610) <= not((layer1_outputs(8859)) xor (layer1_outputs(1198)));
    layer2_outputs(1611) <= not(layer1_outputs(6811)) or (layer1_outputs(9862));
    layer2_outputs(1612) <= (layer1_outputs(7357)) and (layer1_outputs(4185));
    layer2_outputs(1613) <= (layer1_outputs(4947)) and not (layer1_outputs(9659));
    layer2_outputs(1614) <= (layer1_outputs(4747)) and not (layer1_outputs(4283));
    layer2_outputs(1615) <= (layer1_outputs(6863)) and (layer1_outputs(1368));
    layer2_outputs(1616) <= (layer1_outputs(9176)) and not (layer1_outputs(9361));
    layer2_outputs(1617) <= not(layer1_outputs(10057));
    layer2_outputs(1618) <= (layer1_outputs(2883)) or (layer1_outputs(5372));
    layer2_outputs(1619) <= (layer1_outputs(3264)) xor (layer1_outputs(1647));
    layer2_outputs(1620) <= layer1_outputs(557);
    layer2_outputs(1621) <= (layer1_outputs(3416)) and not (layer1_outputs(6528));
    layer2_outputs(1622) <= layer1_outputs(8216);
    layer2_outputs(1623) <= not(layer1_outputs(7641));
    layer2_outputs(1624) <= not((layer1_outputs(3855)) and (layer1_outputs(1152)));
    layer2_outputs(1625) <= not((layer1_outputs(2640)) or (layer1_outputs(1820)));
    layer2_outputs(1626) <= layer1_outputs(7894);
    layer2_outputs(1627) <= layer1_outputs(906);
    layer2_outputs(1628) <= not(layer1_outputs(6956)) or (layer1_outputs(4479));
    layer2_outputs(1629) <= (layer1_outputs(4087)) or (layer1_outputs(5004));
    layer2_outputs(1630) <= not(layer1_outputs(3694));
    layer2_outputs(1631) <= (layer1_outputs(5956)) and (layer1_outputs(9363));
    layer2_outputs(1632) <= not(layer1_outputs(6255)) or (layer1_outputs(1063));
    layer2_outputs(1633) <= layer1_outputs(1649);
    layer2_outputs(1634) <= not(layer1_outputs(5856));
    layer2_outputs(1635) <= not(layer1_outputs(812));
    layer2_outputs(1636) <= not((layer1_outputs(146)) and (layer1_outputs(5535)));
    layer2_outputs(1637) <= not((layer1_outputs(9542)) and (layer1_outputs(8631)));
    layer2_outputs(1638) <= layer1_outputs(3648);
    layer2_outputs(1639) <= (layer1_outputs(3410)) xor (layer1_outputs(4014));
    layer2_outputs(1640) <= not(layer1_outputs(1107));
    layer2_outputs(1641) <= not(layer1_outputs(9099)) or (layer1_outputs(6828));
    layer2_outputs(1642) <= layer1_outputs(6663);
    layer2_outputs(1643) <= not(layer1_outputs(7872));
    layer2_outputs(1644) <= not((layer1_outputs(9159)) or (layer1_outputs(4313)));
    layer2_outputs(1645) <= layer1_outputs(9984);
    layer2_outputs(1646) <= not((layer1_outputs(3256)) and (layer1_outputs(9890)));
    layer2_outputs(1647) <= not(layer1_outputs(9278));
    layer2_outputs(1648) <= (layer1_outputs(2052)) or (layer1_outputs(4949));
    layer2_outputs(1649) <= (layer1_outputs(2907)) xor (layer1_outputs(9447));
    layer2_outputs(1650) <= (layer1_outputs(3098)) and not (layer1_outputs(4058));
    layer2_outputs(1651) <= layer1_outputs(4683);
    layer2_outputs(1652) <= not((layer1_outputs(7668)) or (layer1_outputs(6879)));
    layer2_outputs(1653) <= layer1_outputs(8821);
    layer2_outputs(1654) <= not(layer1_outputs(3693));
    layer2_outputs(1655) <= (layer1_outputs(8666)) and not (layer1_outputs(7349));
    layer2_outputs(1656) <= (layer1_outputs(9105)) and (layer1_outputs(1730));
    layer2_outputs(1657) <= not((layer1_outputs(587)) and (layer1_outputs(620)));
    layer2_outputs(1658) <= (layer1_outputs(5587)) or (layer1_outputs(3341));
    layer2_outputs(1659) <= layer1_outputs(6202);
    layer2_outputs(1660) <= not((layer1_outputs(4388)) and (layer1_outputs(321)));
    layer2_outputs(1661) <= not(layer1_outputs(775));
    layer2_outputs(1662) <= layer1_outputs(8249);
    layer2_outputs(1663) <= layer1_outputs(9756);
    layer2_outputs(1664) <= not((layer1_outputs(6214)) and (layer1_outputs(7959)));
    layer2_outputs(1665) <= not((layer1_outputs(3763)) xor (layer1_outputs(6908)));
    layer2_outputs(1666) <= layer1_outputs(251);
    layer2_outputs(1667) <= (layer1_outputs(8991)) and not (layer1_outputs(5922));
    layer2_outputs(1668) <= layer1_outputs(9788);
    layer2_outputs(1669) <= (layer1_outputs(4870)) xor (layer1_outputs(3830));
    layer2_outputs(1670) <= not(layer1_outputs(9776));
    layer2_outputs(1671) <= not(layer1_outputs(3183)) or (layer1_outputs(1995));
    layer2_outputs(1672) <= not((layer1_outputs(10171)) and (layer1_outputs(7451)));
    layer2_outputs(1673) <= not(layer1_outputs(7309));
    layer2_outputs(1674) <= layer1_outputs(10077);
    layer2_outputs(1675) <= (layer1_outputs(8102)) or (layer1_outputs(9099));
    layer2_outputs(1676) <= not(layer1_outputs(5396));
    layer2_outputs(1677) <= layer1_outputs(8045);
    layer2_outputs(1678) <= (layer1_outputs(3743)) and (layer1_outputs(1179));
    layer2_outputs(1679) <= not((layer1_outputs(6218)) and (layer1_outputs(5827)));
    layer2_outputs(1680) <= (layer1_outputs(2645)) or (layer1_outputs(4185));
    layer2_outputs(1681) <= not((layer1_outputs(8549)) and (layer1_outputs(8807)));
    layer2_outputs(1682) <= layer1_outputs(8237);
    layer2_outputs(1683) <= not((layer1_outputs(5938)) xor (layer1_outputs(10194)));
    layer2_outputs(1684) <= layer1_outputs(9563);
    layer2_outputs(1685) <= not(layer1_outputs(7702));
    layer2_outputs(1686) <= not((layer1_outputs(9933)) xor (layer1_outputs(2741)));
    layer2_outputs(1687) <= not(layer1_outputs(997)) or (layer1_outputs(9504));
    layer2_outputs(1688) <= not(layer1_outputs(3962)) or (layer1_outputs(4126));
    layer2_outputs(1689) <= (layer1_outputs(7782)) and not (layer1_outputs(4776));
    layer2_outputs(1690) <= (layer1_outputs(9303)) or (layer1_outputs(5598));
    layer2_outputs(1691) <= layer1_outputs(1485);
    layer2_outputs(1692) <= (layer1_outputs(5245)) xor (layer1_outputs(3258));
    layer2_outputs(1693) <= (layer1_outputs(9880)) xor (layer1_outputs(8692));
    layer2_outputs(1694) <= layer1_outputs(10159);
    layer2_outputs(1695) <= layer1_outputs(3856);
    layer2_outputs(1696) <= layer1_outputs(1089);
    layer2_outputs(1697) <= not(layer1_outputs(9158));
    layer2_outputs(1698) <= not(layer1_outputs(8486));
    layer2_outputs(1699) <= layer1_outputs(2635);
    layer2_outputs(1700) <= layer1_outputs(6476);
    layer2_outputs(1701) <= not(layer1_outputs(7616));
    layer2_outputs(1702) <= not(layer1_outputs(3639));
    layer2_outputs(1703) <= '1';
    layer2_outputs(1704) <= not((layer1_outputs(8943)) xor (layer1_outputs(9261)));
    layer2_outputs(1705) <= not((layer1_outputs(5646)) and (layer1_outputs(6563)));
    layer2_outputs(1706) <= not(layer1_outputs(4626)) or (layer1_outputs(6838));
    layer2_outputs(1707) <= (layer1_outputs(9949)) xor (layer1_outputs(1130));
    layer2_outputs(1708) <= not(layer1_outputs(324));
    layer2_outputs(1709) <= not(layer1_outputs(8930));
    layer2_outputs(1710) <= layer1_outputs(8171);
    layer2_outputs(1711) <= (layer1_outputs(8432)) xor (layer1_outputs(1593));
    layer2_outputs(1712) <= layer1_outputs(9879);
    layer2_outputs(1713) <= (layer1_outputs(1434)) or (layer1_outputs(10110));
    layer2_outputs(1714) <= (layer1_outputs(996)) and (layer1_outputs(9290));
    layer2_outputs(1715) <= (layer1_outputs(2633)) and not (layer1_outputs(851));
    layer2_outputs(1716) <= layer1_outputs(4539);
    layer2_outputs(1717) <= layer1_outputs(7298);
    layer2_outputs(1718) <= not(layer1_outputs(8586));
    layer2_outputs(1719) <= not(layer1_outputs(10017));
    layer2_outputs(1720) <= (layer1_outputs(1838)) xor (layer1_outputs(9007));
    layer2_outputs(1721) <= layer1_outputs(3807);
    layer2_outputs(1722) <= not((layer1_outputs(9771)) and (layer1_outputs(5682)));
    layer2_outputs(1723) <= not(layer1_outputs(8625));
    layer2_outputs(1724) <= layer1_outputs(2823);
    layer2_outputs(1725) <= layer1_outputs(8069);
    layer2_outputs(1726) <= not(layer1_outputs(7251));
    layer2_outputs(1727) <= not((layer1_outputs(3774)) and (layer1_outputs(3237)));
    layer2_outputs(1728) <= (layer1_outputs(6513)) or (layer1_outputs(1188));
    layer2_outputs(1729) <= not(layer1_outputs(2744)) or (layer1_outputs(7733));
    layer2_outputs(1730) <= (layer1_outputs(3542)) and (layer1_outputs(5613));
    layer2_outputs(1731) <= not(layer1_outputs(4284)) or (layer1_outputs(10135));
    layer2_outputs(1732) <= not(layer1_outputs(5071)) or (layer1_outputs(289));
    layer2_outputs(1733) <= layer1_outputs(4087);
    layer2_outputs(1734) <= layer1_outputs(1346);
    layer2_outputs(1735) <= not(layer1_outputs(9471)) or (layer1_outputs(748));
    layer2_outputs(1736) <= layer1_outputs(9873);
    layer2_outputs(1737) <= not((layer1_outputs(1453)) and (layer1_outputs(1129)));
    layer2_outputs(1738) <= layer1_outputs(8803);
    layer2_outputs(1739) <= (layer1_outputs(3637)) and (layer1_outputs(1397));
    layer2_outputs(1740) <= not(layer1_outputs(3987));
    layer2_outputs(1741) <= layer1_outputs(4954);
    layer2_outputs(1742) <= not(layer1_outputs(507));
    layer2_outputs(1743) <= not((layer1_outputs(8654)) xor (layer1_outputs(4577)));
    layer2_outputs(1744) <= not((layer1_outputs(3462)) or (layer1_outputs(7354)));
    layer2_outputs(1745) <= layer1_outputs(2155);
    layer2_outputs(1746) <= not(layer1_outputs(2269));
    layer2_outputs(1747) <= not((layer1_outputs(1755)) xor (layer1_outputs(1878)));
    layer2_outputs(1748) <= not((layer1_outputs(8265)) xor (layer1_outputs(367)));
    layer2_outputs(1749) <= not(layer1_outputs(1651)) or (layer1_outputs(7665));
    layer2_outputs(1750) <= layer1_outputs(4269);
    layer2_outputs(1751) <= not(layer1_outputs(424));
    layer2_outputs(1752) <= (layer1_outputs(10130)) and (layer1_outputs(8455));
    layer2_outputs(1753) <= not(layer1_outputs(9642));
    layer2_outputs(1754) <= (layer1_outputs(5835)) and not (layer1_outputs(4967));
    layer2_outputs(1755) <= layer1_outputs(9845);
    layer2_outputs(1756) <= not((layer1_outputs(6773)) or (layer1_outputs(2215)));
    layer2_outputs(1757) <= not(layer1_outputs(4732));
    layer2_outputs(1758) <= layer1_outputs(7335);
    layer2_outputs(1759) <= (layer1_outputs(232)) or (layer1_outputs(170));
    layer2_outputs(1760) <= not(layer1_outputs(5667));
    layer2_outputs(1761) <= not(layer1_outputs(4506)) or (layer1_outputs(3824));
    layer2_outputs(1762) <= not((layer1_outputs(7047)) xor (layer1_outputs(5244)));
    layer2_outputs(1763) <= (layer1_outputs(1591)) and not (layer1_outputs(8708));
    layer2_outputs(1764) <= not(layer1_outputs(2481)) or (layer1_outputs(5833));
    layer2_outputs(1765) <= layer1_outputs(4919);
    layer2_outputs(1766) <= not(layer1_outputs(6495));
    layer2_outputs(1767) <= layer1_outputs(8246);
    layer2_outputs(1768) <= layer1_outputs(9548);
    layer2_outputs(1769) <= not((layer1_outputs(1208)) or (layer1_outputs(5227)));
    layer2_outputs(1770) <= not(layer1_outputs(3466)) or (layer1_outputs(283));
    layer2_outputs(1771) <= not(layer1_outputs(5820));
    layer2_outputs(1772) <= not((layer1_outputs(3147)) xor (layer1_outputs(3558)));
    layer2_outputs(1773) <= not(layer1_outputs(1940)) or (layer1_outputs(7032));
    layer2_outputs(1774) <= not(layer1_outputs(9037));
    layer2_outputs(1775) <= not((layer1_outputs(3701)) or (layer1_outputs(4737)));
    layer2_outputs(1776) <= (layer1_outputs(8186)) xor (layer1_outputs(8549));
    layer2_outputs(1777) <= not(layer1_outputs(873)) or (layer1_outputs(9501));
    layer2_outputs(1778) <= layer1_outputs(6390);
    layer2_outputs(1779) <= not(layer1_outputs(9332));
    layer2_outputs(1780) <= (layer1_outputs(204)) and (layer1_outputs(4813));
    layer2_outputs(1781) <= layer1_outputs(10023);
    layer2_outputs(1782) <= layer1_outputs(9055);
    layer2_outputs(1783) <= not((layer1_outputs(630)) and (layer1_outputs(3496)));
    layer2_outputs(1784) <= layer1_outputs(4054);
    layer2_outputs(1785) <= layer1_outputs(7529);
    layer2_outputs(1786) <= not((layer1_outputs(2353)) and (layer1_outputs(5112)));
    layer2_outputs(1787) <= not(layer1_outputs(3287));
    layer2_outputs(1788) <= not((layer1_outputs(4174)) and (layer1_outputs(1741)));
    layer2_outputs(1789) <= not(layer1_outputs(634)) or (layer1_outputs(931));
    layer2_outputs(1790) <= not((layer1_outputs(3966)) xor (layer1_outputs(3227)));
    layer2_outputs(1791) <= not(layer1_outputs(1471)) or (layer1_outputs(2528));
    layer2_outputs(1792) <= not(layer1_outputs(753));
    layer2_outputs(1793) <= layer1_outputs(4971);
    layer2_outputs(1794) <= not(layer1_outputs(888));
    layer2_outputs(1795) <= not(layer1_outputs(1221));
    layer2_outputs(1796) <= layer1_outputs(4537);
    layer2_outputs(1797) <= not(layer1_outputs(572)) or (layer1_outputs(9429));
    layer2_outputs(1798) <= layer1_outputs(6919);
    layer2_outputs(1799) <= not(layer1_outputs(8457));
    layer2_outputs(1800) <= not((layer1_outputs(595)) xor (layer1_outputs(5325)));
    layer2_outputs(1801) <= not(layer1_outputs(640));
    layer2_outputs(1802) <= (layer1_outputs(1360)) xor (layer1_outputs(3615));
    layer2_outputs(1803) <= not(layer1_outputs(9939));
    layer2_outputs(1804) <= (layer1_outputs(751)) and (layer1_outputs(994));
    layer2_outputs(1805) <= layer1_outputs(6806);
    layer2_outputs(1806) <= not(layer1_outputs(9498));
    layer2_outputs(1807) <= layer1_outputs(6158);
    layer2_outputs(1808) <= layer1_outputs(330);
    layer2_outputs(1809) <= (layer1_outputs(4001)) or (layer1_outputs(5766));
    layer2_outputs(1810) <= not((layer1_outputs(4800)) and (layer1_outputs(3735)));
    layer2_outputs(1811) <= layer1_outputs(6629);
    layer2_outputs(1812) <= layer1_outputs(5042);
    layer2_outputs(1813) <= not((layer1_outputs(9731)) and (layer1_outputs(3747)));
    layer2_outputs(1814) <= not((layer1_outputs(302)) and (layer1_outputs(938)));
    layer2_outputs(1815) <= (layer1_outputs(2152)) and not (layer1_outputs(7557));
    layer2_outputs(1816) <= layer1_outputs(7709);
    layer2_outputs(1817) <= (layer1_outputs(8156)) xor (layer1_outputs(3518));
    layer2_outputs(1818) <= not(layer1_outputs(6422));
    layer2_outputs(1819) <= layer1_outputs(1284);
    layer2_outputs(1820) <= not((layer1_outputs(156)) or (layer1_outputs(4449)));
    layer2_outputs(1821) <= not(layer1_outputs(3469)) or (layer1_outputs(3182));
    layer2_outputs(1822) <= '0';
    layer2_outputs(1823) <= (layer1_outputs(9265)) and not (layer1_outputs(10128));
    layer2_outputs(1824) <= not((layer1_outputs(8851)) and (layer1_outputs(10164)));
    layer2_outputs(1825) <= not((layer1_outputs(9549)) and (layer1_outputs(9977)));
    layer2_outputs(1826) <= not(layer1_outputs(8231)) or (layer1_outputs(3707));
    layer2_outputs(1827) <= not((layer1_outputs(99)) or (layer1_outputs(3439)));
    layer2_outputs(1828) <= '0';
    layer2_outputs(1829) <= not(layer1_outputs(963));
    layer2_outputs(1830) <= '0';
    layer2_outputs(1831) <= layer1_outputs(1560);
    layer2_outputs(1832) <= layer1_outputs(7191);
    layer2_outputs(1833) <= not(layer1_outputs(1739));
    layer2_outputs(1834) <= (layer1_outputs(9969)) and (layer1_outputs(4488));
    layer2_outputs(1835) <= layer1_outputs(6520);
    layer2_outputs(1836) <= not(layer1_outputs(8939)) or (layer1_outputs(4291));
    layer2_outputs(1837) <= (layer1_outputs(4221)) and not (layer1_outputs(6605));
    layer2_outputs(1838) <= layer1_outputs(7631);
    layer2_outputs(1839) <= layer1_outputs(5715);
    layer2_outputs(1840) <= not((layer1_outputs(9475)) xor (layer1_outputs(7995)));
    layer2_outputs(1841) <= layer1_outputs(7727);
    layer2_outputs(1842) <= (layer1_outputs(10048)) or (layer1_outputs(4579));
    layer2_outputs(1843) <= layer1_outputs(4183);
    layer2_outputs(1844) <= (layer1_outputs(6855)) xor (layer1_outputs(5578));
    layer2_outputs(1845) <= not(layer1_outputs(699));
    layer2_outputs(1846) <= (layer1_outputs(1318)) xor (layer1_outputs(9188));
    layer2_outputs(1847) <= not(layer1_outputs(6701)) or (layer1_outputs(6998));
    layer2_outputs(1848) <= (layer1_outputs(3799)) and not (layer1_outputs(2748));
    layer2_outputs(1849) <= not((layer1_outputs(8157)) or (layer1_outputs(8956)));
    layer2_outputs(1850) <= layer1_outputs(2372);
    layer2_outputs(1851) <= not((layer1_outputs(8885)) and (layer1_outputs(10072)));
    layer2_outputs(1852) <= not(layer1_outputs(5488));
    layer2_outputs(1853) <= (layer1_outputs(1096)) and not (layer1_outputs(5158));
    layer2_outputs(1854) <= '0';
    layer2_outputs(1855) <= not(layer1_outputs(4952));
    layer2_outputs(1856) <= not(layer1_outputs(4526));
    layer2_outputs(1857) <= (layer1_outputs(9779)) and not (layer1_outputs(2532));
    layer2_outputs(1858) <= (layer1_outputs(9986)) or (layer1_outputs(3886));
    layer2_outputs(1859) <= not(layer1_outputs(4336));
    layer2_outputs(1860) <= '0';
    layer2_outputs(1861) <= layer1_outputs(4810);
    layer2_outputs(1862) <= not((layer1_outputs(9947)) or (layer1_outputs(9263)));
    layer2_outputs(1863) <= (layer1_outputs(2166)) and not (layer1_outputs(166));
    layer2_outputs(1864) <= (layer1_outputs(1333)) and (layer1_outputs(3481));
    layer2_outputs(1865) <= layer1_outputs(6834);
    layer2_outputs(1866) <= not(layer1_outputs(7515));
    layer2_outputs(1867) <= not((layer1_outputs(2089)) or (layer1_outputs(829)));
    layer2_outputs(1868) <= not((layer1_outputs(2796)) and (layer1_outputs(608)));
    layer2_outputs(1869) <= not(layer1_outputs(4021));
    layer2_outputs(1870) <= (layer1_outputs(4173)) and not (layer1_outputs(1991));
    layer2_outputs(1871) <= not((layer1_outputs(4196)) xor (layer1_outputs(4459)));
    layer2_outputs(1872) <= not((layer1_outputs(5462)) xor (layer1_outputs(4431)));
    layer2_outputs(1873) <= layer1_outputs(2327);
    layer2_outputs(1874) <= not(layer1_outputs(10161));
    layer2_outputs(1875) <= (layer1_outputs(6630)) xor (layer1_outputs(170));
    layer2_outputs(1876) <= not(layer1_outputs(5548)) or (layer1_outputs(2615));
    layer2_outputs(1877) <= not(layer1_outputs(5716)) or (layer1_outputs(1323));
    layer2_outputs(1878) <= not(layer1_outputs(2165));
    layer2_outputs(1879) <= (layer1_outputs(2622)) xor (layer1_outputs(5986));
    layer2_outputs(1880) <= (layer1_outputs(226)) and not (layer1_outputs(3634));
    layer2_outputs(1881) <= not(layer1_outputs(9287));
    layer2_outputs(1882) <= not(layer1_outputs(2199));
    layer2_outputs(1883) <= layer1_outputs(10019);
    layer2_outputs(1884) <= (layer1_outputs(6791)) xor (layer1_outputs(7565));
    layer2_outputs(1885) <= (layer1_outputs(10012)) and not (layer1_outputs(1957));
    layer2_outputs(1886) <= not(layer1_outputs(1768));
    layer2_outputs(1887) <= not(layer1_outputs(5932)) or (layer1_outputs(9481));
    layer2_outputs(1888) <= (layer1_outputs(5976)) and not (layer1_outputs(7169));
    layer2_outputs(1889) <= not(layer1_outputs(3678)) or (layer1_outputs(6778));
    layer2_outputs(1890) <= not((layer1_outputs(8719)) xor (layer1_outputs(7867)));
    layer2_outputs(1891) <= layer1_outputs(8740);
    layer2_outputs(1892) <= layer1_outputs(9360);
    layer2_outputs(1893) <= (layer1_outputs(6425)) and not (layer1_outputs(2884));
    layer2_outputs(1894) <= layer1_outputs(4271);
    layer2_outputs(1895) <= (layer1_outputs(6089)) and not (layer1_outputs(5725));
    layer2_outputs(1896) <= not(layer1_outputs(5094));
    layer2_outputs(1897) <= layer1_outputs(6065);
    layer2_outputs(1898) <= not((layer1_outputs(8932)) and (layer1_outputs(6141)));
    layer2_outputs(1899) <= layer1_outputs(9641);
    layer2_outputs(1900) <= not(layer1_outputs(5016));
    layer2_outputs(1901) <= not(layer1_outputs(5368)) or (layer1_outputs(7743));
    layer2_outputs(1902) <= (layer1_outputs(6962)) xor (layer1_outputs(2453));
    layer2_outputs(1903) <= not(layer1_outputs(7217)) or (layer1_outputs(10020));
    layer2_outputs(1904) <= (layer1_outputs(8865)) and not (layer1_outputs(3170));
    layer2_outputs(1905) <= layer1_outputs(432);
    layer2_outputs(1906) <= layer1_outputs(3624);
    layer2_outputs(1907) <= (layer1_outputs(2674)) and not (layer1_outputs(7372));
    layer2_outputs(1908) <= not(layer1_outputs(6627)) or (layer1_outputs(672));
    layer2_outputs(1909) <= not(layer1_outputs(522));
    layer2_outputs(1910) <= layer1_outputs(516);
    layer2_outputs(1911) <= (layer1_outputs(7834)) and not (layer1_outputs(7622));
    layer2_outputs(1912) <= not(layer1_outputs(834));
    layer2_outputs(1913) <= (layer1_outputs(2781)) or (layer1_outputs(6721));
    layer2_outputs(1914) <= not(layer1_outputs(6735));
    layer2_outputs(1915) <= layer1_outputs(8971);
    layer2_outputs(1916) <= not(layer1_outputs(2907));
    layer2_outputs(1917) <= not(layer1_outputs(7497));
    layer2_outputs(1918) <= layer1_outputs(10036);
    layer2_outputs(1919) <= '1';
    layer2_outputs(1920) <= not(layer1_outputs(5651));
    layer2_outputs(1921) <= (layer1_outputs(1402)) xor (layer1_outputs(476));
    layer2_outputs(1922) <= layer1_outputs(2762);
    layer2_outputs(1923) <= layer1_outputs(2381);
    layer2_outputs(1924) <= layer1_outputs(7254);
    layer2_outputs(1925) <= layer1_outputs(9689);
    layer2_outputs(1926) <= not((layer1_outputs(1168)) xor (layer1_outputs(1706)));
    layer2_outputs(1927) <= layer1_outputs(3912);
    layer2_outputs(1928) <= (layer1_outputs(1186)) and (layer1_outputs(3463));
    layer2_outputs(1929) <= (layer1_outputs(6071)) and not (layer1_outputs(10154));
    layer2_outputs(1930) <= not(layer1_outputs(5683));
    layer2_outputs(1931) <= not((layer1_outputs(4122)) and (layer1_outputs(5424)));
    layer2_outputs(1932) <= not(layer1_outputs(2464));
    layer2_outputs(1933) <= not(layer1_outputs(370)) or (layer1_outputs(8751));
    layer2_outputs(1934) <= not(layer1_outputs(1705));
    layer2_outputs(1935) <= not(layer1_outputs(7280)) or (layer1_outputs(4426));
    layer2_outputs(1936) <= not((layer1_outputs(5172)) xor (layer1_outputs(8824)));
    layer2_outputs(1937) <= (layer1_outputs(4769)) or (layer1_outputs(5866));
    layer2_outputs(1938) <= (layer1_outputs(9594)) and not (layer1_outputs(9648));
    layer2_outputs(1939) <= not((layer1_outputs(2205)) xor (layer1_outputs(1327)));
    layer2_outputs(1940) <= not(layer1_outputs(2442)) or (layer1_outputs(4721));
    layer2_outputs(1941) <= not(layer1_outputs(9208)) or (layer1_outputs(3234));
    layer2_outputs(1942) <= (layer1_outputs(2523)) xor (layer1_outputs(5170));
    layer2_outputs(1943) <= (layer1_outputs(490)) and not (layer1_outputs(10035));
    layer2_outputs(1944) <= not(layer1_outputs(7502)) or (layer1_outputs(740));
    layer2_outputs(1945) <= not(layer1_outputs(5037));
    layer2_outputs(1946) <= (layer1_outputs(9264)) and not (layer1_outputs(6288));
    layer2_outputs(1947) <= not(layer1_outputs(3456));
    layer2_outputs(1948) <= not(layer1_outputs(9181));
    layer2_outputs(1949) <= (layer1_outputs(2614)) or (layer1_outputs(1783));
    layer2_outputs(1950) <= (layer1_outputs(8315)) or (layer1_outputs(7153));
    layer2_outputs(1951) <= (layer1_outputs(7323)) or (layer1_outputs(8678));
    layer2_outputs(1952) <= layer1_outputs(2666);
    layer2_outputs(1953) <= layer1_outputs(7421);
    layer2_outputs(1954) <= not(layer1_outputs(5825)) or (layer1_outputs(9848));
    layer2_outputs(1955) <= (layer1_outputs(2637)) or (layer1_outputs(8411));
    layer2_outputs(1956) <= not(layer1_outputs(9629));
    layer2_outputs(1957) <= (layer1_outputs(6501)) xor (layer1_outputs(7522));
    layer2_outputs(1958) <= not(layer1_outputs(7345));
    layer2_outputs(1959) <= layer1_outputs(1816);
    layer2_outputs(1960) <= not(layer1_outputs(1849)) or (layer1_outputs(9493));
    layer2_outputs(1961) <= layer1_outputs(8027);
    layer2_outputs(1962) <= layer1_outputs(414);
    layer2_outputs(1963) <= not(layer1_outputs(6429));
    layer2_outputs(1964) <= layer1_outputs(5562);
    layer2_outputs(1965) <= not(layer1_outputs(1868));
    layer2_outputs(1966) <= (layer1_outputs(10028)) and (layer1_outputs(6800));
    layer2_outputs(1967) <= not(layer1_outputs(897));
    layer2_outputs(1968) <= (layer1_outputs(2694)) xor (layer1_outputs(6820));
    layer2_outputs(1969) <= not(layer1_outputs(200)) or (layer1_outputs(6160));
    layer2_outputs(1970) <= not((layer1_outputs(830)) or (layer1_outputs(9252)));
    layer2_outputs(1971) <= layer1_outputs(5634);
    layer2_outputs(1972) <= (layer1_outputs(7819)) and (layer1_outputs(6306));
    layer2_outputs(1973) <= layer1_outputs(934);
    layer2_outputs(1974) <= (layer1_outputs(6029)) and (layer1_outputs(7585));
    layer2_outputs(1975) <= layer1_outputs(7238);
    layer2_outputs(1976) <= layer1_outputs(4627);
    layer2_outputs(1977) <= not(layer1_outputs(7577));
    layer2_outputs(1978) <= not((layer1_outputs(1117)) or (layer1_outputs(1047)));
    layer2_outputs(1979) <= not(layer1_outputs(7075));
    layer2_outputs(1980) <= layer1_outputs(9595);
    layer2_outputs(1981) <= layer1_outputs(4740);
    layer2_outputs(1982) <= not(layer1_outputs(9296));
    layer2_outputs(1983) <= layer1_outputs(5776);
    layer2_outputs(1984) <= not((layer1_outputs(9918)) and (layer1_outputs(6805)));
    layer2_outputs(1985) <= not((layer1_outputs(3181)) xor (layer1_outputs(1646)));
    layer2_outputs(1986) <= layer1_outputs(970);
    layer2_outputs(1987) <= not(layer1_outputs(6170));
    layer2_outputs(1988) <= not(layer1_outputs(8150));
    layer2_outputs(1989) <= not(layer1_outputs(4474));
    layer2_outputs(1990) <= not(layer1_outputs(9296));
    layer2_outputs(1991) <= layer1_outputs(9179);
    layer2_outputs(1992) <= not((layer1_outputs(529)) and (layer1_outputs(9625)));
    layer2_outputs(1993) <= not(layer1_outputs(8970));
    layer2_outputs(1994) <= (layer1_outputs(2041)) and not (layer1_outputs(4065));
    layer2_outputs(1995) <= not((layer1_outputs(6360)) and (layer1_outputs(2377)));
    layer2_outputs(1996) <= '1';
    layer2_outputs(1997) <= not(layer1_outputs(5426));
    layer2_outputs(1998) <= not(layer1_outputs(1409));
    layer2_outputs(1999) <= not(layer1_outputs(912));
    layer2_outputs(2000) <= not(layer1_outputs(6416));
    layer2_outputs(2001) <= layer1_outputs(5285);
    layer2_outputs(2002) <= (layer1_outputs(9392)) and (layer1_outputs(10005));
    layer2_outputs(2003) <= not((layer1_outputs(1711)) xor (layer1_outputs(2923)));
    layer2_outputs(2004) <= not((layer1_outputs(3238)) or (layer1_outputs(9079)));
    layer2_outputs(2005) <= not(layer1_outputs(7633));
    layer2_outputs(2006) <= not(layer1_outputs(7394));
    layer2_outputs(2007) <= layer1_outputs(3);
    layer2_outputs(2008) <= not(layer1_outputs(6868));
    layer2_outputs(2009) <= (layer1_outputs(10200)) and not (layer1_outputs(1713));
    layer2_outputs(2010) <= layer1_outputs(6581);
    layer2_outputs(2011) <= not((layer1_outputs(1477)) and (layer1_outputs(4969)));
    layer2_outputs(2012) <= layer1_outputs(5243);
    layer2_outputs(2013) <= (layer1_outputs(4836)) xor (layer1_outputs(8609));
    layer2_outputs(2014) <= not(layer1_outputs(7564));
    layer2_outputs(2015) <= layer1_outputs(4238);
    layer2_outputs(2016) <= not(layer1_outputs(7866));
    layer2_outputs(2017) <= not(layer1_outputs(4772));
    layer2_outputs(2018) <= not((layer1_outputs(7909)) or (layer1_outputs(8442)));
    layer2_outputs(2019) <= layer1_outputs(1394);
    layer2_outputs(2020) <= not(layer1_outputs(10158));
    layer2_outputs(2021) <= not((layer1_outputs(3274)) xor (layer1_outputs(8524)));
    layer2_outputs(2022) <= layer1_outputs(4716);
    layer2_outputs(2023) <= layer1_outputs(2063);
    layer2_outputs(2024) <= not((layer1_outputs(8850)) or (layer1_outputs(3574)));
    layer2_outputs(2025) <= not(layer1_outputs(5914)) or (layer1_outputs(4998));
    layer2_outputs(2026) <= layer1_outputs(10016);
    layer2_outputs(2027) <= not(layer1_outputs(8183)) or (layer1_outputs(9457));
    layer2_outputs(2028) <= (layer1_outputs(3671)) and (layer1_outputs(3853));
    layer2_outputs(2029) <= layer1_outputs(1922);
    layer2_outputs(2030) <= layer1_outputs(7418);
    layer2_outputs(2031) <= not(layer1_outputs(1187));
    layer2_outputs(2032) <= (layer1_outputs(1252)) and not (layer1_outputs(126));
    layer2_outputs(2033) <= layer1_outputs(69);
    layer2_outputs(2034) <= (layer1_outputs(2543)) and (layer1_outputs(9395));
    layer2_outputs(2035) <= '0';
    layer2_outputs(2036) <= not((layer1_outputs(1929)) or (layer1_outputs(1141)));
    layer2_outputs(2037) <= (layer1_outputs(5176)) and not (layer1_outputs(8681));
    layer2_outputs(2038) <= layer1_outputs(7507);
    layer2_outputs(2039) <= not((layer1_outputs(1070)) and (layer1_outputs(9221)));
    layer2_outputs(2040) <= (layer1_outputs(565)) or (layer1_outputs(6536));
    layer2_outputs(2041) <= not(layer1_outputs(3210));
    layer2_outputs(2042) <= not((layer1_outputs(8481)) and (layer1_outputs(7413)));
    layer2_outputs(2043) <= (layer1_outputs(4570)) and not (layer1_outputs(9131));
    layer2_outputs(2044) <= not(layer1_outputs(3552));
    layer2_outputs(2045) <= not((layer1_outputs(5810)) and (layer1_outputs(9463)));
    layer2_outputs(2046) <= (layer1_outputs(4308)) or (layer1_outputs(5147));
    layer2_outputs(2047) <= not((layer1_outputs(2371)) and (layer1_outputs(4658)));
    layer2_outputs(2048) <= not(layer1_outputs(606));
    layer2_outputs(2049) <= (layer1_outputs(2963)) xor (layer1_outputs(6969));
    layer2_outputs(2050) <= layer1_outputs(9786);
    layer2_outputs(2051) <= (layer1_outputs(5195)) and not (layer1_outputs(3995));
    layer2_outputs(2052) <= not(layer1_outputs(7674)) or (layer1_outputs(2310));
    layer2_outputs(2053) <= layer1_outputs(2521);
    layer2_outputs(2054) <= not(layer1_outputs(4158)) or (layer1_outputs(4261));
    layer2_outputs(2055) <= not(layer1_outputs(4599)) or (layer1_outputs(1298));
    layer2_outputs(2056) <= not(layer1_outputs(3066));
    layer2_outputs(2057) <= (layer1_outputs(1733)) and not (layer1_outputs(3636));
    layer2_outputs(2058) <= (layer1_outputs(6104)) xor (layer1_outputs(1907));
    layer2_outputs(2059) <= not((layer1_outputs(4899)) and (layer1_outputs(309)));
    layer2_outputs(2060) <= layer1_outputs(3348);
    layer2_outputs(2061) <= not((layer1_outputs(5485)) xor (layer1_outputs(1764)));
    layer2_outputs(2062) <= not(layer1_outputs(9372)) or (layer1_outputs(4759));
    layer2_outputs(2063) <= not(layer1_outputs(3798)) or (layer1_outputs(5884));
    layer2_outputs(2064) <= layer1_outputs(9660);
    layer2_outputs(2065) <= (layer1_outputs(6257)) or (layer1_outputs(847));
    layer2_outputs(2066) <= (layer1_outputs(1142)) xor (layer1_outputs(5618));
    layer2_outputs(2067) <= not((layer1_outputs(9533)) and (layer1_outputs(3580)));
    layer2_outputs(2068) <= layer1_outputs(4175);
    layer2_outputs(2069) <= layer1_outputs(3377);
    layer2_outputs(2070) <= not(layer1_outputs(6297));
    layer2_outputs(2071) <= (layer1_outputs(3498)) and not (layer1_outputs(7103));
    layer2_outputs(2072) <= not(layer1_outputs(10120));
    layer2_outputs(2073) <= layer1_outputs(6318);
    layer2_outputs(2074) <= not(layer1_outputs(10177));
    layer2_outputs(2075) <= layer1_outputs(6684);
    layer2_outputs(2076) <= not(layer1_outputs(8881));
    layer2_outputs(2077) <= (layer1_outputs(4562)) and not (layer1_outputs(6413));
    layer2_outputs(2078) <= not(layer1_outputs(6902));
    layer2_outputs(2079) <= (layer1_outputs(2909)) and not (layer1_outputs(9546));
    layer2_outputs(2080) <= layer1_outputs(6125);
    layer2_outputs(2081) <= not(layer1_outputs(7964));
    layer2_outputs(2082) <= (layer1_outputs(1375)) or (layer1_outputs(1712));
    layer2_outputs(2083) <= (layer1_outputs(377)) and not (layer1_outputs(3534));
    layer2_outputs(2084) <= not(layer1_outputs(7661));
    layer2_outputs(2085) <= (layer1_outputs(6862)) or (layer1_outputs(7472));
    layer2_outputs(2086) <= not((layer1_outputs(8275)) xor (layer1_outputs(6034)));
    layer2_outputs(2087) <= not(layer1_outputs(8420)) or (layer1_outputs(2039));
    layer2_outputs(2088) <= (layer1_outputs(7400)) and (layer1_outputs(1253));
    layer2_outputs(2089) <= not(layer1_outputs(9028));
    layer2_outputs(2090) <= layer1_outputs(2484);
    layer2_outputs(2091) <= not(layer1_outputs(4007));
    layer2_outputs(2092) <= (layer1_outputs(2114)) and (layer1_outputs(7009));
    layer2_outputs(2093) <= not(layer1_outputs(10208));
    layer2_outputs(2094) <= not(layer1_outputs(5185));
    layer2_outputs(2095) <= (layer1_outputs(4134)) and not (layer1_outputs(2836));
    layer2_outputs(2096) <= layer1_outputs(2193);
    layer2_outputs(2097) <= (layer1_outputs(1457)) and not (layer1_outputs(4452));
    layer2_outputs(2098) <= not(layer1_outputs(6421));
    layer2_outputs(2099) <= layer1_outputs(3640);
    layer2_outputs(2100) <= layer1_outputs(4392);
    layer2_outputs(2101) <= not(layer1_outputs(5177)) or (layer1_outputs(9257));
    layer2_outputs(2102) <= not(layer1_outputs(2012)) or (layer1_outputs(4922));
    layer2_outputs(2103) <= not(layer1_outputs(1866));
    layer2_outputs(2104) <= not(layer1_outputs(7796)) or (layer1_outputs(7919));
    layer2_outputs(2105) <= not(layer1_outputs(2803));
    layer2_outputs(2106) <= not(layer1_outputs(4596)) or (layer1_outputs(2870));
    layer2_outputs(2107) <= (layer1_outputs(3081)) and not (layer1_outputs(1899));
    layer2_outputs(2108) <= (layer1_outputs(8180)) or (layer1_outputs(2065));
    layer2_outputs(2109) <= not(layer1_outputs(1696));
    layer2_outputs(2110) <= not((layer1_outputs(9717)) or (layer1_outputs(2828)));
    layer2_outputs(2111) <= layer1_outputs(6092);
    layer2_outputs(2112) <= (layer1_outputs(4251)) or (layer1_outputs(8767));
    layer2_outputs(2113) <= layer1_outputs(1412);
    layer2_outputs(2114) <= layer1_outputs(7987);
    layer2_outputs(2115) <= not((layer1_outputs(6243)) xor (layer1_outputs(10094)));
    layer2_outputs(2116) <= layer1_outputs(9734);
    layer2_outputs(2117) <= not((layer1_outputs(3942)) xor (layer1_outputs(9930)));
    layer2_outputs(2118) <= not(layer1_outputs(3498)) or (layer1_outputs(7940));
    layer2_outputs(2119) <= layer1_outputs(6427);
    layer2_outputs(2120) <= (layer1_outputs(7481)) and (layer1_outputs(799));
    layer2_outputs(2121) <= '0';
    layer2_outputs(2122) <= layer1_outputs(1692);
    layer2_outputs(2123) <= not((layer1_outputs(7216)) and (layer1_outputs(1888)));
    layer2_outputs(2124) <= layer1_outputs(2174);
    layer2_outputs(2125) <= not(layer1_outputs(4505));
    layer2_outputs(2126) <= not(layer1_outputs(3355)) or (layer1_outputs(57));
    layer2_outputs(2127) <= (layer1_outputs(6164)) and not (layer1_outputs(6961));
    layer2_outputs(2128) <= layer1_outputs(4944);
    layer2_outputs(2129) <= not(layer1_outputs(787)) or (layer1_outputs(483));
    layer2_outputs(2130) <= (layer1_outputs(6397)) and (layer1_outputs(6173));
    layer2_outputs(2131) <= not(layer1_outputs(1471)) or (layer1_outputs(2369));
    layer2_outputs(2132) <= (layer1_outputs(302)) and (layer1_outputs(1947));
    layer2_outputs(2133) <= not(layer1_outputs(6253));
    layer2_outputs(2134) <= layer1_outputs(7838);
    layer2_outputs(2135) <= layer1_outputs(8704);
    layer2_outputs(2136) <= layer1_outputs(1582);
    layer2_outputs(2137) <= not(layer1_outputs(2564));
    layer2_outputs(2138) <= not((layer1_outputs(7073)) or (layer1_outputs(651)));
    layer2_outputs(2139) <= (layer1_outputs(4436)) or (layer1_outputs(1354));
    layer2_outputs(2140) <= not(layer1_outputs(4794));
    layer2_outputs(2141) <= not((layer1_outputs(8275)) and (layer1_outputs(5110)));
    layer2_outputs(2142) <= not(layer1_outputs(3413)) or (layer1_outputs(4392));
    layer2_outputs(2143) <= not(layer1_outputs(7016)) or (layer1_outputs(7754));
    layer2_outputs(2144) <= not(layer1_outputs(8259));
    layer2_outputs(2145) <= not(layer1_outputs(5006)) or (layer1_outputs(7886));
    layer2_outputs(2146) <= not(layer1_outputs(9321));
    layer2_outputs(2147) <= (layer1_outputs(6770)) xor (layer1_outputs(10130));
    layer2_outputs(2148) <= layer1_outputs(3680);
    layer2_outputs(2149) <= (layer1_outputs(9462)) and not (layer1_outputs(4620));
    layer2_outputs(2150) <= layer1_outputs(8270);
    layer2_outputs(2151) <= layer1_outputs(9058);
    layer2_outputs(2152) <= (layer1_outputs(1039)) and not (layer1_outputs(2571));
    layer2_outputs(2153) <= not(layer1_outputs(6523));
    layer2_outputs(2154) <= (layer1_outputs(5385)) xor (layer1_outputs(10042));
    layer2_outputs(2155) <= not(layer1_outputs(1087));
    layer2_outputs(2156) <= not(layer1_outputs(5172));
    layer2_outputs(2157) <= '0';
    layer2_outputs(2158) <= layer1_outputs(1322);
    layer2_outputs(2159) <= '1';
    layer2_outputs(2160) <= not(layer1_outputs(7511));
    layer2_outputs(2161) <= layer1_outputs(6136);
    layer2_outputs(2162) <= layer1_outputs(6789);
    layer2_outputs(2163) <= not(layer1_outputs(6239));
    layer2_outputs(2164) <= not(layer1_outputs(2445));
    layer2_outputs(2165) <= not(layer1_outputs(4611));
    layer2_outputs(2166) <= layer1_outputs(3225);
    layer2_outputs(2167) <= '0';
    layer2_outputs(2168) <= (layer1_outputs(1856)) xor (layer1_outputs(8052));
    layer2_outputs(2169) <= not(layer1_outputs(9478));
    layer2_outputs(2170) <= (layer1_outputs(4753)) and (layer1_outputs(402));
    layer2_outputs(2171) <= layer1_outputs(8116);
    layer2_outputs(2172) <= not((layer1_outputs(6696)) or (layer1_outputs(4334)));
    layer2_outputs(2173) <= not((layer1_outputs(3184)) and (layer1_outputs(7501)));
    layer2_outputs(2174) <= layer1_outputs(3629);
    layer2_outputs(2175) <= not((layer1_outputs(5142)) xor (layer1_outputs(5612)));
    layer2_outputs(2176) <= (layer1_outputs(1396)) xor (layer1_outputs(3751));
    layer2_outputs(2177) <= layer1_outputs(6881);
    layer2_outputs(2178) <= (layer1_outputs(8533)) xor (layer1_outputs(9100));
    layer2_outputs(2179) <= layer1_outputs(6248);
    layer2_outputs(2180) <= not((layer1_outputs(7891)) or (layer1_outputs(4403)));
    layer2_outputs(2181) <= not(layer1_outputs(5207)) or (layer1_outputs(1634));
    layer2_outputs(2182) <= (layer1_outputs(2684)) and not (layer1_outputs(9390));
    layer2_outputs(2183) <= not((layer1_outputs(776)) xor (layer1_outputs(3795)));
    layer2_outputs(2184) <= not(layer1_outputs(9475)) or (layer1_outputs(2159));
    layer2_outputs(2185) <= '0';
    layer2_outputs(2186) <= not(layer1_outputs(8021)) or (layer1_outputs(1239));
    layer2_outputs(2187) <= not(layer1_outputs(1350));
    layer2_outputs(2188) <= not((layer1_outputs(2529)) or (layer1_outputs(5606)));
    layer2_outputs(2189) <= (layer1_outputs(7863)) or (layer1_outputs(3958));
    layer2_outputs(2190) <= layer1_outputs(9057);
    layer2_outputs(2191) <= not((layer1_outputs(2964)) xor (layer1_outputs(4595)));
    layer2_outputs(2192) <= not((layer1_outputs(6814)) xor (layer1_outputs(7596)));
    layer2_outputs(2193) <= layer1_outputs(7745);
    layer2_outputs(2194) <= not(layer1_outputs(8706)) or (layer1_outputs(6303));
    layer2_outputs(2195) <= layer1_outputs(6737);
    layer2_outputs(2196) <= layer1_outputs(4189);
    layer2_outputs(2197) <= not(layer1_outputs(6484));
    layer2_outputs(2198) <= (layer1_outputs(5976)) and not (layer1_outputs(2962));
    layer2_outputs(2199) <= layer1_outputs(4959);
    layer2_outputs(2200) <= (layer1_outputs(9938)) xor (layer1_outputs(6592));
    layer2_outputs(2201) <= layer1_outputs(9266);
    layer2_outputs(2202) <= layer1_outputs(3380);
    layer2_outputs(2203) <= not(layer1_outputs(8799)) or (layer1_outputs(2393));
    layer2_outputs(2204) <= not((layer1_outputs(4225)) xor (layer1_outputs(7110)));
    layer2_outputs(2205) <= not(layer1_outputs(1220));
    layer2_outputs(2206) <= layer1_outputs(4513);
    layer2_outputs(2207) <= not(layer1_outputs(9487));
    layer2_outputs(2208) <= not((layer1_outputs(9016)) xor (layer1_outputs(8170)));
    layer2_outputs(2209) <= layer1_outputs(3532);
    layer2_outputs(2210) <= not((layer1_outputs(6607)) and (layer1_outputs(4875)));
    layer2_outputs(2211) <= (layer1_outputs(1289)) and not (layer1_outputs(7112));
    layer2_outputs(2212) <= not(layer1_outputs(3443));
    layer2_outputs(2213) <= not((layer1_outputs(9337)) and (layer1_outputs(3541)));
    layer2_outputs(2214) <= (layer1_outputs(5321)) or (layer1_outputs(6670));
    layer2_outputs(2215) <= not(layer1_outputs(9612));
    layer2_outputs(2216) <= not(layer1_outputs(3871));
    layer2_outputs(2217) <= (layer1_outputs(6485)) and (layer1_outputs(7349));
    layer2_outputs(2218) <= layer1_outputs(3072);
    layer2_outputs(2219) <= not(layer1_outputs(6956)) or (layer1_outputs(8482));
    layer2_outputs(2220) <= layer1_outputs(718);
    layer2_outputs(2221) <= not(layer1_outputs(7424)) or (layer1_outputs(4317));
    layer2_outputs(2222) <= not(layer1_outputs(536));
    layer2_outputs(2223) <= (layer1_outputs(1514)) and not (layer1_outputs(6143));
    layer2_outputs(2224) <= not(layer1_outputs(9791));
    layer2_outputs(2225) <= not(layer1_outputs(9123)) or (layer1_outputs(8334));
    layer2_outputs(2226) <= not(layer1_outputs(891));
    layer2_outputs(2227) <= (layer1_outputs(10191)) and not (layer1_outputs(6490));
    layer2_outputs(2228) <= layer1_outputs(2772);
    layer2_outputs(2229) <= not(layer1_outputs(5425)) or (layer1_outputs(2870));
    layer2_outputs(2230) <= not(layer1_outputs(798)) or (layer1_outputs(1663));
    layer2_outputs(2231) <= not((layer1_outputs(280)) and (layer1_outputs(4204)));
    layer2_outputs(2232) <= not(layer1_outputs(8518));
    layer2_outputs(2233) <= (layer1_outputs(8543)) and not (layer1_outputs(9013));
    layer2_outputs(2234) <= not(layer1_outputs(7179)) or (layer1_outputs(6026));
    layer2_outputs(2235) <= (layer1_outputs(3478)) xor (layer1_outputs(7464));
    layer2_outputs(2236) <= (layer1_outputs(2760)) and (layer1_outputs(4902));
    layer2_outputs(2237) <= (layer1_outputs(9112)) and (layer1_outputs(3374));
    layer2_outputs(2238) <= layer1_outputs(7301);
    layer2_outputs(2239) <= not(layer1_outputs(8308));
    layer2_outputs(2240) <= not((layer1_outputs(3585)) xor (layer1_outputs(504)));
    layer2_outputs(2241) <= not(layer1_outputs(3132));
    layer2_outputs(2242) <= not(layer1_outputs(3314));
    layer2_outputs(2243) <= layer1_outputs(8556);
    layer2_outputs(2244) <= not((layer1_outputs(941)) xor (layer1_outputs(2267)));
    layer2_outputs(2245) <= not(layer1_outputs(4908));
    layer2_outputs(2246) <= (layer1_outputs(3246)) or (layer1_outputs(192));
    layer2_outputs(2247) <= (layer1_outputs(9733)) xor (layer1_outputs(1182));
    layer2_outputs(2248) <= layer1_outputs(2317);
    layer2_outputs(2249) <= layer1_outputs(880);
    layer2_outputs(2250) <= not(layer1_outputs(2528));
    layer2_outputs(2251) <= (layer1_outputs(9388)) xor (layer1_outputs(9142));
    layer2_outputs(2252) <= not((layer1_outputs(1525)) xor (layer1_outputs(7341)));
    layer2_outputs(2253) <= layer1_outputs(4088);
    layer2_outputs(2254) <= not((layer1_outputs(8713)) or (layer1_outputs(6017)));
    layer2_outputs(2255) <= not((layer1_outputs(3152)) or (layer1_outputs(1492)));
    layer2_outputs(2256) <= not(layer1_outputs(3710));
    layer2_outputs(2257) <= (layer1_outputs(2499)) and not (layer1_outputs(1464));
    layer2_outputs(2258) <= not((layer1_outputs(5983)) xor (layer1_outputs(5032)));
    layer2_outputs(2259) <= not(layer1_outputs(1705)) or (layer1_outputs(4070));
    layer2_outputs(2260) <= (layer1_outputs(8075)) and not (layer1_outputs(3157));
    layer2_outputs(2261) <= layer1_outputs(5406);
    layer2_outputs(2262) <= not(layer1_outputs(6112)) or (layer1_outputs(953));
    layer2_outputs(2263) <= not((layer1_outputs(4375)) or (layer1_outputs(2644)));
    layer2_outputs(2264) <= not(layer1_outputs(8916));
    layer2_outputs(2265) <= not((layer1_outputs(5415)) or (layer1_outputs(3784)));
    layer2_outputs(2266) <= layer1_outputs(9893);
    layer2_outputs(2267) <= (layer1_outputs(5741)) xor (layer1_outputs(220));
    layer2_outputs(2268) <= (layer1_outputs(5330)) and not (layer1_outputs(6011));
    layer2_outputs(2269) <= layer1_outputs(535);
    layer2_outputs(2270) <= not(layer1_outputs(3037));
    layer2_outputs(2271) <= (layer1_outputs(7411)) or (layer1_outputs(4845));
    layer2_outputs(2272) <= layer1_outputs(5109);
    layer2_outputs(2273) <= (layer1_outputs(2236)) xor (layer1_outputs(1154));
    layer2_outputs(2274) <= not((layer1_outputs(9359)) and (layer1_outputs(6453)));
    layer2_outputs(2275) <= (layer1_outputs(7688)) and not (layer1_outputs(5332));
    layer2_outputs(2276) <= layer1_outputs(3501);
    layer2_outputs(2277) <= layer1_outputs(3137);
    layer2_outputs(2278) <= (layer1_outputs(2779)) xor (layer1_outputs(9973));
    layer2_outputs(2279) <= not(layer1_outputs(5967)) or (layer1_outputs(5403));
    layer2_outputs(2280) <= layer1_outputs(205);
    layer2_outputs(2281) <= not((layer1_outputs(4351)) xor (layer1_outputs(4544)));
    layer2_outputs(2282) <= not((layer1_outputs(9802)) or (layer1_outputs(10101)));
    layer2_outputs(2283) <= layer1_outputs(771);
    layer2_outputs(2284) <= not((layer1_outputs(6764)) or (layer1_outputs(3986)));
    layer2_outputs(2285) <= (layer1_outputs(133)) and (layer1_outputs(3817));
    layer2_outputs(2286) <= not(layer1_outputs(7909));
    layer2_outputs(2287) <= (layer1_outputs(971)) and (layer1_outputs(7503));
    layer2_outputs(2288) <= (layer1_outputs(4619)) and (layer1_outputs(5448));
    layer2_outputs(2289) <= not(layer1_outputs(5498));
    layer2_outputs(2290) <= not(layer1_outputs(7259)) or (layer1_outputs(5423));
    layer2_outputs(2291) <= (layer1_outputs(7684)) and not (layer1_outputs(1602));
    layer2_outputs(2292) <= layer1_outputs(4280);
    layer2_outputs(2293) <= not(layer1_outputs(5818));
    layer2_outputs(2294) <= not(layer1_outputs(4448));
    layer2_outputs(2295) <= not(layer1_outputs(519)) or (layer1_outputs(5057));
    layer2_outputs(2296) <= layer1_outputs(7786);
    layer2_outputs(2297) <= not(layer1_outputs(5933)) or (layer1_outputs(4422));
    layer2_outputs(2298) <= layer1_outputs(6803);
    layer2_outputs(2299) <= not(layer1_outputs(1146));
    layer2_outputs(2300) <= (layer1_outputs(1920)) or (layer1_outputs(3923));
    layer2_outputs(2301) <= not(layer1_outputs(6038));
    layer2_outputs(2302) <= (layer1_outputs(9031)) or (layer1_outputs(9288));
    layer2_outputs(2303) <= (layer1_outputs(371)) or (layer1_outputs(1659));
    layer2_outputs(2304) <= layer1_outputs(8676);
    layer2_outputs(2305) <= not(layer1_outputs(5270));
    layer2_outputs(2306) <= not(layer1_outputs(6731));
    layer2_outputs(2307) <= (layer1_outputs(1138)) xor (layer1_outputs(3308));
    layer2_outputs(2308) <= (layer1_outputs(3833)) and (layer1_outputs(10006));
    layer2_outputs(2309) <= not(layer1_outputs(5580)) or (layer1_outputs(8967));
    layer2_outputs(2310) <= not(layer1_outputs(5560));
    layer2_outputs(2311) <= layer1_outputs(5720);
    layer2_outputs(2312) <= layer1_outputs(1675);
    layer2_outputs(2313) <= not((layer1_outputs(7336)) xor (layer1_outputs(482)));
    layer2_outputs(2314) <= not(layer1_outputs(1994));
    layer2_outputs(2315) <= (layer1_outputs(5601)) xor (layer1_outputs(8290));
    layer2_outputs(2316) <= (layer1_outputs(6221)) and not (layer1_outputs(9031));
    layer2_outputs(2317) <= layer1_outputs(3608);
    layer2_outputs(2318) <= not((layer1_outputs(8947)) xor (layer1_outputs(1197)));
    layer2_outputs(2319) <= (layer1_outputs(5281)) and (layer1_outputs(2521));
    layer2_outputs(2320) <= not(layer1_outputs(859)) or (layer1_outputs(6891));
    layer2_outputs(2321) <= (layer1_outputs(1515)) and not (layer1_outputs(8964));
    layer2_outputs(2322) <= not((layer1_outputs(7734)) xor (layer1_outputs(8415)));
    layer2_outputs(2323) <= layer1_outputs(7564);
    layer2_outputs(2324) <= layer1_outputs(3633);
    layer2_outputs(2325) <= not(layer1_outputs(4685));
    layer2_outputs(2326) <= (layer1_outputs(8534)) xor (layer1_outputs(4150));
    layer2_outputs(2327) <= (layer1_outputs(2745)) and not (layer1_outputs(2707));
    layer2_outputs(2328) <= not(layer1_outputs(2687)) or (layer1_outputs(4354));
    layer2_outputs(2329) <= not((layer1_outputs(8812)) and (layer1_outputs(9649)));
    layer2_outputs(2330) <= layer1_outputs(7390);
    layer2_outputs(2331) <= (layer1_outputs(4474)) and not (layer1_outputs(3866));
    layer2_outputs(2332) <= not(layer1_outputs(9657));
    layer2_outputs(2333) <= layer1_outputs(638);
    layer2_outputs(2334) <= not((layer1_outputs(7730)) xor (layer1_outputs(3384)));
    layer2_outputs(2335) <= not(layer1_outputs(2210)) or (layer1_outputs(5210));
    layer2_outputs(2336) <= not(layer1_outputs(3336));
    layer2_outputs(2337) <= '0';
    layer2_outputs(2338) <= not(layer1_outputs(4606));
    layer2_outputs(2339) <= (layer1_outputs(1461)) or (layer1_outputs(5249));
    layer2_outputs(2340) <= not(layer1_outputs(2700)) or (layer1_outputs(3890));
    layer2_outputs(2341) <= (layer1_outputs(9777)) and not (layer1_outputs(229));
    layer2_outputs(2342) <= layer1_outputs(3509);
    layer2_outputs(2343) <= (layer1_outputs(5395)) and (layer1_outputs(8047));
    layer2_outputs(2344) <= layer1_outputs(5547);
    layer2_outputs(2345) <= layer1_outputs(6600);
    layer2_outputs(2346) <= layer1_outputs(158);
    layer2_outputs(2347) <= layer1_outputs(8691);
    layer2_outputs(2348) <= not((layer1_outputs(9205)) xor (layer1_outputs(8490)));
    layer2_outputs(2349) <= layer1_outputs(6827);
    layer2_outputs(2350) <= not(layer1_outputs(5514)) or (layer1_outputs(2407));
    layer2_outputs(2351) <= (layer1_outputs(3423)) and (layer1_outputs(1154));
    layer2_outputs(2352) <= not(layer1_outputs(5320));
    layer2_outputs(2353) <= not(layer1_outputs(9572)) or (layer1_outputs(8205));
    layer2_outputs(2354) <= (layer1_outputs(6295)) and not (layer1_outputs(666));
    layer2_outputs(2355) <= layer1_outputs(346);
    layer2_outputs(2356) <= layer1_outputs(4680);
    layer2_outputs(2357) <= layer1_outputs(8596);
    layer2_outputs(2358) <= not(layer1_outputs(4904));
    layer2_outputs(2359) <= (layer1_outputs(9139)) xor (layer1_outputs(7610));
    layer2_outputs(2360) <= (layer1_outputs(2840)) and (layer1_outputs(6958));
    layer2_outputs(2361) <= layer1_outputs(510);
    layer2_outputs(2362) <= '1';
    layer2_outputs(2363) <= not((layer1_outputs(6762)) xor (layer1_outputs(6583)));
    layer2_outputs(2364) <= (layer1_outputs(6036)) and not (layer1_outputs(9120));
    layer2_outputs(2365) <= (layer1_outputs(9333)) or (layer1_outputs(9374));
    layer2_outputs(2366) <= not(layer1_outputs(4510));
    layer2_outputs(2367) <= (layer1_outputs(9698)) or (layer1_outputs(3550));
    layer2_outputs(2368) <= (layer1_outputs(5664)) xor (layer1_outputs(6361));
    layer2_outputs(2369) <= not(layer1_outputs(1691));
    layer2_outputs(2370) <= not(layer1_outputs(4710));
    layer2_outputs(2371) <= not((layer1_outputs(2373)) xor (layer1_outputs(34)));
    layer2_outputs(2372) <= not(layer1_outputs(6222));
    layer2_outputs(2373) <= not(layer1_outputs(5739)) or (layer1_outputs(7643));
    layer2_outputs(2374) <= not(layer1_outputs(6349));
    layer2_outputs(2375) <= not(layer1_outputs(2356));
    layer2_outputs(2376) <= not(layer1_outputs(1525));
    layer2_outputs(2377) <= (layer1_outputs(2742)) or (layer1_outputs(4372));
    layer2_outputs(2378) <= layer1_outputs(5506);
    layer2_outputs(2379) <= (layer1_outputs(2859)) xor (layer1_outputs(5023));
    layer2_outputs(2380) <= layer1_outputs(5869);
    layer2_outputs(2381) <= not((layer1_outputs(7119)) or (layer1_outputs(3690)));
    layer2_outputs(2382) <= not((layer1_outputs(7865)) xor (layer1_outputs(1426)));
    layer2_outputs(2383) <= layer1_outputs(4369);
    layer2_outputs(2384) <= layer1_outputs(10180);
    layer2_outputs(2385) <= layer1_outputs(2431);
    layer2_outputs(2386) <= layer1_outputs(5706);
    layer2_outputs(2387) <= not((layer1_outputs(5322)) xor (layer1_outputs(1949)));
    layer2_outputs(2388) <= not((layer1_outputs(3495)) or (layer1_outputs(4141)));
    layer2_outputs(2389) <= not(layer1_outputs(8446));
    layer2_outputs(2390) <= layer1_outputs(4426);
    layer2_outputs(2391) <= not((layer1_outputs(7825)) xor (layer1_outputs(10203)));
    layer2_outputs(2392) <= layer1_outputs(477);
    layer2_outputs(2393) <= not(layer1_outputs(6552));
    layer2_outputs(2394) <= layer1_outputs(4149);
    layer2_outputs(2395) <= not(layer1_outputs(3688));
    layer2_outputs(2396) <= layer1_outputs(3318);
    layer2_outputs(2397) <= not(layer1_outputs(450));
    layer2_outputs(2398) <= not(layer1_outputs(659));
    layer2_outputs(2399) <= layer1_outputs(7507);
    layer2_outputs(2400) <= not(layer1_outputs(2059));
    layer2_outputs(2401) <= '1';
    layer2_outputs(2402) <= (layer1_outputs(6653)) or (layer1_outputs(9941));
    layer2_outputs(2403) <= not(layer1_outputs(8180));
    layer2_outputs(2404) <= not(layer1_outputs(2626));
    layer2_outputs(2405) <= not(layer1_outputs(2760)) or (layer1_outputs(6379));
    layer2_outputs(2406) <= layer1_outputs(6048);
    layer2_outputs(2407) <= (layer1_outputs(6152)) xor (layer1_outputs(2578));
    layer2_outputs(2408) <= not(layer1_outputs(1058));
    layer2_outputs(2409) <= not(layer1_outputs(5723));
    layer2_outputs(2410) <= not((layer1_outputs(10213)) or (layer1_outputs(1593)));
    layer2_outputs(2411) <= not(layer1_outputs(3428));
    layer2_outputs(2412) <= not(layer1_outputs(6548)) or (layer1_outputs(9609));
    layer2_outputs(2413) <= not(layer1_outputs(314)) or (layer1_outputs(4206));
    layer2_outputs(2414) <= (layer1_outputs(9515)) xor (layer1_outputs(5431));
    layer2_outputs(2415) <= layer1_outputs(8977);
    layer2_outputs(2416) <= not(layer1_outputs(7855));
    layer2_outputs(2417) <= (layer1_outputs(7039)) or (layer1_outputs(6518));
    layer2_outputs(2418) <= layer1_outputs(5963);
    layer2_outputs(2419) <= not(layer1_outputs(1544));
    layer2_outputs(2420) <= not(layer1_outputs(9515));
    layer2_outputs(2421) <= not((layer1_outputs(2443)) or (layer1_outputs(9098)));
    layer2_outputs(2422) <= not(layer1_outputs(5717)) or (layer1_outputs(6171));
    layer2_outputs(2423) <= not((layer1_outputs(988)) xor (layer1_outputs(2270)));
    layer2_outputs(2424) <= (layer1_outputs(9615)) or (layer1_outputs(1714));
    layer2_outputs(2425) <= (layer1_outputs(64)) and not (layer1_outputs(2988));
    layer2_outputs(2426) <= layer1_outputs(4446);
    layer2_outputs(2427) <= (layer1_outputs(10086)) xor (layer1_outputs(3128));
    layer2_outputs(2428) <= not(layer1_outputs(2660));
    layer2_outputs(2429) <= layer1_outputs(483);
    layer2_outputs(2430) <= not(layer1_outputs(1878));
    layer2_outputs(2431) <= not(layer1_outputs(8255));
    layer2_outputs(2432) <= not(layer1_outputs(537));
    layer2_outputs(2433) <= layer1_outputs(3659);
    layer2_outputs(2434) <= layer1_outputs(8978);
    layer2_outputs(2435) <= (layer1_outputs(470)) or (layer1_outputs(2987));
    layer2_outputs(2436) <= (layer1_outputs(9508)) xor (layer1_outputs(7659));
    layer2_outputs(2437) <= (layer1_outputs(7544)) or (layer1_outputs(1668));
    layer2_outputs(2438) <= layer1_outputs(6196);
    layer2_outputs(2439) <= not(layer1_outputs(6904)) or (layer1_outputs(802));
    layer2_outputs(2440) <= not((layer1_outputs(5805)) and (layer1_outputs(1011)));
    layer2_outputs(2441) <= not(layer1_outputs(7795));
    layer2_outputs(2442) <= layer1_outputs(2687);
    layer2_outputs(2443) <= layer1_outputs(9072);
    layer2_outputs(2444) <= (layer1_outputs(2715)) and not (layer1_outputs(1963));
    layer2_outputs(2445) <= not(layer1_outputs(5984));
    layer2_outputs(2446) <= layer1_outputs(3708);
    layer2_outputs(2447) <= not((layer1_outputs(4176)) and (layer1_outputs(3461)));
    layer2_outputs(2448) <= (layer1_outputs(4843)) and (layer1_outputs(4035));
    layer2_outputs(2449) <= (layer1_outputs(1299)) and (layer1_outputs(8864));
    layer2_outputs(2450) <= layer1_outputs(6157);
    layer2_outputs(2451) <= '1';
    layer2_outputs(2452) <= not(layer1_outputs(148)) or (layer1_outputs(8623));
    layer2_outputs(2453) <= layer1_outputs(8580);
    layer2_outputs(2454) <= layer1_outputs(9012);
    layer2_outputs(2455) <= not((layer1_outputs(5898)) xor (layer1_outputs(8758)));
    layer2_outputs(2456) <= layer1_outputs(2945);
    layer2_outputs(2457) <= layer1_outputs(3671);
    layer2_outputs(2458) <= not(layer1_outputs(2359));
    layer2_outputs(2459) <= (layer1_outputs(2969)) or (layer1_outputs(3769));
    layer2_outputs(2460) <= (layer1_outputs(2772)) and (layer1_outputs(2030));
    layer2_outputs(2461) <= layer1_outputs(197);
    layer2_outputs(2462) <= (layer1_outputs(7678)) or (layer1_outputs(6412));
    layer2_outputs(2463) <= layer1_outputs(2222);
    layer2_outputs(2464) <= not(layer1_outputs(8295)) or (layer1_outputs(2264));
    layer2_outputs(2465) <= (layer1_outputs(5397)) and (layer1_outputs(1041));
    layer2_outputs(2466) <= not((layer1_outputs(6076)) or (layer1_outputs(5532)));
    layer2_outputs(2467) <= layer1_outputs(6111);
    layer2_outputs(2468) <= (layer1_outputs(8421)) and (layer1_outputs(9224));
    layer2_outputs(2469) <= (layer1_outputs(1713)) xor (layer1_outputs(8817));
    layer2_outputs(2470) <= not((layer1_outputs(7731)) or (layer1_outputs(5568)));
    layer2_outputs(2471) <= not(layer1_outputs(3637));
    layer2_outputs(2472) <= layer1_outputs(8344);
    layer2_outputs(2473) <= not(layer1_outputs(2428)) or (layer1_outputs(6930));
    layer2_outputs(2474) <= not(layer1_outputs(5828));
    layer2_outputs(2475) <= layer1_outputs(4441);
    layer2_outputs(2476) <= layer1_outputs(1077);
    layer2_outputs(2477) <= layer1_outputs(6681);
    layer2_outputs(2478) <= not((layer1_outputs(5711)) or (layer1_outputs(3178)));
    layer2_outputs(2479) <= not(layer1_outputs(8438));
    layer2_outputs(2480) <= not((layer1_outputs(5300)) xor (layer1_outputs(2581)));
    layer2_outputs(2481) <= (layer1_outputs(6912)) and not (layer1_outputs(7723));
    layer2_outputs(2482) <= (layer1_outputs(9713)) and (layer1_outputs(1279));
    layer2_outputs(2483) <= not((layer1_outputs(3963)) xor (layer1_outputs(6345)));
    layer2_outputs(2484) <= (layer1_outputs(1113)) and not (layer1_outputs(1364));
    layer2_outputs(2485) <= not((layer1_outputs(4495)) xor (layer1_outputs(6777)));
    layer2_outputs(2486) <= not((layer1_outputs(1623)) or (layer1_outputs(2955)));
    layer2_outputs(2487) <= (layer1_outputs(864)) or (layer1_outputs(189));
    layer2_outputs(2488) <= not(layer1_outputs(9526)) or (layer1_outputs(3121));
    layer2_outputs(2489) <= not(layer1_outputs(7707)) or (layer1_outputs(6293));
    layer2_outputs(2490) <= not(layer1_outputs(7775));
    layer2_outputs(2491) <= not(layer1_outputs(2351));
    layer2_outputs(2492) <= layer1_outputs(9304);
    layer2_outputs(2493) <= layer1_outputs(3101);
    layer2_outputs(2494) <= layer1_outputs(2701);
    layer2_outputs(2495) <= (layer1_outputs(7770)) and not (layer1_outputs(6068));
    layer2_outputs(2496) <= layer1_outputs(5851);
    layer2_outputs(2497) <= layer1_outputs(5062);
    layer2_outputs(2498) <= not(layer1_outputs(3310));
    layer2_outputs(2499) <= not(layer1_outputs(6926)) or (layer1_outputs(8676));
    layer2_outputs(2500) <= not(layer1_outputs(4494));
    layer2_outputs(2501) <= (layer1_outputs(10021)) xor (layer1_outputs(3864));
    layer2_outputs(2502) <= not((layer1_outputs(6950)) or (layer1_outputs(3960)));
    layer2_outputs(2503) <= not(layer1_outputs(8272));
    layer2_outputs(2504) <= (layer1_outputs(1003)) xor (layer1_outputs(9905));
    layer2_outputs(2505) <= (layer1_outputs(8243)) and not (layer1_outputs(3213));
    layer2_outputs(2506) <= not((layer1_outputs(8559)) and (layer1_outputs(2305)));
    layer2_outputs(2507) <= not(layer1_outputs(2607));
    layer2_outputs(2508) <= (layer1_outputs(3098)) and not (layer1_outputs(6003));
    layer2_outputs(2509) <= layer1_outputs(7682);
    layer2_outputs(2510) <= (layer1_outputs(9267)) and not (layer1_outputs(5440));
    layer2_outputs(2511) <= (layer1_outputs(4953)) and not (layer1_outputs(6988));
    layer2_outputs(2512) <= (layer1_outputs(5855)) and not (layer1_outputs(5296));
    layer2_outputs(2513) <= (layer1_outputs(9953)) and not (layer1_outputs(9580));
    layer2_outputs(2514) <= (layer1_outputs(4987)) and not (layer1_outputs(8878));
    layer2_outputs(2515) <= (layer1_outputs(9931)) xor (layer1_outputs(1556));
    layer2_outputs(2516) <= not(layer1_outputs(6108));
    layer2_outputs(2517) <= layer1_outputs(2253);
    layer2_outputs(2518) <= not(layer1_outputs(1941)) or (layer1_outputs(1571));
    layer2_outputs(2519) <= (layer1_outputs(658)) and not (layer1_outputs(2558));
    layer2_outputs(2520) <= not((layer1_outputs(430)) xor (layer1_outputs(3529)));
    layer2_outputs(2521) <= (layer1_outputs(6717)) xor (layer1_outputs(4981));
    layer2_outputs(2522) <= (layer1_outputs(3356)) and not (layer1_outputs(4767));
    layer2_outputs(2523) <= layer1_outputs(168);
    layer2_outputs(2524) <= not(layer1_outputs(9255));
    layer2_outputs(2525) <= (layer1_outputs(9757)) and (layer1_outputs(2559));
    layer2_outputs(2526) <= not(layer1_outputs(1279));
    layer2_outputs(2527) <= not(layer1_outputs(199));
    layer2_outputs(2528) <= layer1_outputs(342);
    layer2_outputs(2529) <= '0';
    layer2_outputs(2530) <= layer1_outputs(8343);
    layer2_outputs(2531) <= (layer1_outputs(340)) xor (layer1_outputs(5439));
    layer2_outputs(2532) <= not((layer1_outputs(502)) xor (layer1_outputs(2886)));
    layer2_outputs(2533) <= layer1_outputs(8337);
    layer2_outputs(2534) <= layer1_outputs(6015);
    layer2_outputs(2535) <= (layer1_outputs(2537)) or (layer1_outputs(9928));
    layer2_outputs(2536) <= (layer1_outputs(6687)) and not (layer1_outputs(8339));
    layer2_outputs(2537) <= layer1_outputs(1473);
    layer2_outputs(2538) <= not(layer1_outputs(3471));
    layer2_outputs(2539) <= not((layer1_outputs(9483)) or (layer1_outputs(3073)));
    layer2_outputs(2540) <= not(layer1_outputs(5643)) or (layer1_outputs(7854));
    layer2_outputs(2541) <= not(layer1_outputs(4668)) or (layer1_outputs(6418));
    layer2_outputs(2542) <= (layer1_outputs(8230)) or (layer1_outputs(1130));
    layer2_outputs(2543) <= not(layer1_outputs(5760));
    layer2_outputs(2544) <= layer1_outputs(5593);
    layer2_outputs(2545) <= layer1_outputs(7271);
    layer2_outputs(2546) <= not(layer1_outputs(6135));
    layer2_outputs(2547) <= (layer1_outputs(2075)) and not (layer1_outputs(6925));
    layer2_outputs(2548) <= not(layer1_outputs(5317)) or (layer1_outputs(2900));
    layer2_outputs(2549) <= (layer1_outputs(2582)) and not (layer1_outputs(4927));
    layer2_outputs(2550) <= not(layer1_outputs(3400));
    layer2_outputs(2551) <= not((layer1_outputs(9973)) or (layer1_outputs(6778)));
    layer2_outputs(2552) <= not((layer1_outputs(6675)) or (layer1_outputs(7577)));
    layer2_outputs(2553) <= (layer1_outputs(2820)) or (layer1_outputs(2324));
    layer2_outputs(2554) <= not(layer1_outputs(2692));
    layer2_outputs(2555) <= (layer1_outputs(9108)) and not (layer1_outputs(7999));
    layer2_outputs(2556) <= not((layer1_outputs(2045)) and (layer1_outputs(5237)));
    layer2_outputs(2557) <= not(layer1_outputs(4991));
    layer2_outputs(2558) <= layer1_outputs(2299);
    layer2_outputs(2559) <= not((layer1_outputs(3686)) xor (layer1_outputs(5510)));
    layer2_outputs(2560) <= not(layer1_outputs(7023));
    layer2_outputs(2561) <= not(layer1_outputs(3172));
    layer2_outputs(2562) <= (layer1_outputs(9506)) and not (layer1_outputs(4055));
    layer2_outputs(2563) <= layer1_outputs(5232);
    layer2_outputs(2564) <= not(layer1_outputs(4413));
    layer2_outputs(2565) <= '0';
    layer2_outputs(2566) <= (layer1_outputs(1254)) and not (layer1_outputs(3467));
    layer2_outputs(2567) <= layer1_outputs(1770);
    layer2_outputs(2568) <= not((layer1_outputs(1892)) xor (layer1_outputs(3766)));
    layer2_outputs(2569) <= not(layer1_outputs(7983));
    layer2_outputs(2570) <= not((layer1_outputs(7008)) xor (layer1_outputs(9085)));
    layer2_outputs(2571) <= not(layer1_outputs(3876));
    layer2_outputs(2572) <= (layer1_outputs(2736)) and (layer1_outputs(7479));
    layer2_outputs(2573) <= not(layer1_outputs(3929)) or (layer1_outputs(1189));
    layer2_outputs(2574) <= layer1_outputs(9579);
    layer2_outputs(2575) <= (layer1_outputs(2191)) xor (layer1_outputs(7489));
    layer2_outputs(2576) <= not(layer1_outputs(4405));
    layer2_outputs(2577) <= not(layer1_outputs(6121));
    layer2_outputs(2578) <= not(layer1_outputs(9579));
    layer2_outputs(2579) <= (layer1_outputs(2416)) and (layer1_outputs(7205));
    layer2_outputs(2580) <= layer1_outputs(10076);
    layer2_outputs(2581) <= not(layer1_outputs(9798));
    layer2_outputs(2582) <= not(layer1_outputs(9009));
    layer2_outputs(2583) <= layer1_outputs(7883);
    layer2_outputs(2584) <= layer1_outputs(2554);
    layer2_outputs(2585) <= layer1_outputs(3086);
    layer2_outputs(2586) <= not((layer1_outputs(5357)) xor (layer1_outputs(10052)));
    layer2_outputs(2587) <= (layer1_outputs(6129)) xor (layer1_outputs(2096));
    layer2_outputs(2588) <= '0';
    layer2_outputs(2589) <= not((layer1_outputs(9993)) xor (layer1_outputs(2261)));
    layer2_outputs(2590) <= not(layer1_outputs(9116));
    layer2_outputs(2591) <= not(layer1_outputs(2144));
    layer2_outputs(2592) <= not((layer1_outputs(9537)) and (layer1_outputs(9313)));
    layer2_outputs(2593) <= layer1_outputs(320);
    layer2_outputs(2594) <= (layer1_outputs(3240)) xor (layer1_outputs(3306));
    layer2_outputs(2595) <= layer1_outputs(5997);
    layer2_outputs(2596) <= layer1_outputs(6259);
    layer2_outputs(2597) <= (layer1_outputs(4159)) and (layer1_outputs(198));
    layer2_outputs(2598) <= layer1_outputs(3530);
    layer2_outputs(2599) <= layer1_outputs(810);
    layer2_outputs(2600) <= not(layer1_outputs(554));
    layer2_outputs(2601) <= (layer1_outputs(698)) or (layer1_outputs(4982));
    layer2_outputs(2602) <= not(layer1_outputs(2277));
    layer2_outputs(2603) <= layer1_outputs(7288);
    layer2_outputs(2604) <= not(layer1_outputs(5459));
    layer2_outputs(2605) <= (layer1_outputs(1007)) and not (layer1_outputs(2947));
    layer2_outputs(2606) <= not(layer1_outputs(2574));
    layer2_outputs(2607) <= not(layer1_outputs(10065)) or (layer1_outputs(4417));
    layer2_outputs(2608) <= (layer1_outputs(197)) and (layer1_outputs(4521));
    layer2_outputs(2609) <= not(layer1_outputs(9449)) or (layer1_outputs(3704));
    layer2_outputs(2610) <= (layer1_outputs(5554)) or (layer1_outputs(8579));
    layer2_outputs(2611) <= '0';
    layer2_outputs(2612) <= not(layer1_outputs(3562));
    layer2_outputs(2613) <= layer1_outputs(533);
    layer2_outputs(2614) <= not((layer1_outputs(8399)) and (layer1_outputs(7531)));
    layer2_outputs(2615) <= layer1_outputs(1761);
    layer2_outputs(2616) <= layer1_outputs(6080);
    layer2_outputs(2617) <= not(layer1_outputs(3262));
    layer2_outputs(2618) <= (layer1_outputs(5320)) and not (layer1_outputs(9049));
    layer2_outputs(2619) <= not(layer1_outputs(5457));
    layer2_outputs(2620) <= (layer1_outputs(53)) and not (layer1_outputs(7087));
    layer2_outputs(2621) <= not(layer1_outputs(622));
    layer2_outputs(2622) <= not(layer1_outputs(1047));
    layer2_outputs(2623) <= (layer1_outputs(5424)) xor (layer1_outputs(5412));
    layer2_outputs(2624) <= not((layer1_outputs(585)) and (layer1_outputs(9259)));
    layer2_outputs(2625) <= (layer1_outputs(609)) and not (layer1_outputs(7133));
    layer2_outputs(2626) <= layer1_outputs(9914);
    layer2_outputs(2627) <= (layer1_outputs(2332)) xor (layer1_outputs(7625));
    layer2_outputs(2628) <= (layer1_outputs(1934)) xor (layer1_outputs(6833));
    layer2_outputs(2629) <= layer1_outputs(2973);
    layer2_outputs(2630) <= layer1_outputs(309);
    layer2_outputs(2631) <= not(layer1_outputs(2057)) or (layer1_outputs(5022));
    layer2_outputs(2632) <= (layer1_outputs(4093)) and not (layer1_outputs(2715));
    layer2_outputs(2633) <= not(layer1_outputs(2406));
    layer2_outputs(2634) <= layer1_outputs(9669);
    layer2_outputs(2635) <= layer1_outputs(2496);
    layer2_outputs(2636) <= not(layer1_outputs(9654)) or (layer1_outputs(7360));
    layer2_outputs(2637) <= (layer1_outputs(5257)) and not (layer1_outputs(4826));
    layer2_outputs(2638) <= not(layer1_outputs(8592));
    layer2_outputs(2639) <= layer1_outputs(4301);
    layer2_outputs(2640) <= '1';
    layer2_outputs(2641) <= layer1_outputs(86);
    layer2_outputs(2642) <= not(layer1_outputs(897));
    layer2_outputs(2643) <= not((layer1_outputs(2342)) or (layer1_outputs(2837)));
    layer2_outputs(2644) <= not(layer1_outputs(1384));
    layer2_outputs(2645) <= (layer1_outputs(998)) or (layer1_outputs(6399));
    layer2_outputs(2646) <= (layer1_outputs(7468)) xor (layer1_outputs(461));
    layer2_outputs(2647) <= (layer1_outputs(9977)) xor (layer1_outputs(9216));
    layer2_outputs(2648) <= not(layer1_outputs(6058));
    layer2_outputs(2649) <= layer1_outputs(8260);
    layer2_outputs(2650) <= not((layer1_outputs(6936)) xor (layer1_outputs(277)));
    layer2_outputs(2651) <= (layer1_outputs(984)) xor (layer1_outputs(3668));
    layer2_outputs(2652) <= layer1_outputs(1676);
    layer2_outputs(2653) <= not(layer1_outputs(6477));
    layer2_outputs(2654) <= not((layer1_outputs(796)) or (layer1_outputs(9773)));
    layer2_outputs(2655) <= not(layer1_outputs(2525));
    layer2_outputs(2656) <= not(layer1_outputs(7872));
    layer2_outputs(2657) <= (layer1_outputs(10038)) xor (layer1_outputs(2095));
    layer2_outputs(2658) <= layer1_outputs(768);
    layer2_outputs(2659) <= not(layer1_outputs(5895));
    layer2_outputs(2660) <= (layer1_outputs(8812)) and (layer1_outputs(6705));
    layer2_outputs(2661) <= not(layer1_outputs(1056)) or (layer1_outputs(7767));
    layer2_outputs(2662) <= layer1_outputs(4255);
    layer2_outputs(2663) <= '0';
    layer2_outputs(2664) <= layer1_outputs(289);
    layer2_outputs(2665) <= not((layer1_outputs(7429)) xor (layer1_outputs(9958)));
    layer2_outputs(2666) <= (layer1_outputs(3370)) and not (layer1_outputs(7623));
    layer2_outputs(2667) <= layer1_outputs(2507);
    layer2_outputs(2668) <= (layer1_outputs(2318)) and (layer1_outputs(3945));
    layer2_outputs(2669) <= not(layer1_outputs(6109));
    layer2_outputs(2670) <= not(layer1_outputs(8449));
    layer2_outputs(2671) <= not(layer1_outputs(1494));
    layer2_outputs(2672) <= layer1_outputs(4758);
    layer2_outputs(2673) <= layer1_outputs(534);
    layer2_outputs(2674) <= not((layer1_outputs(8083)) and (layer1_outputs(6546)));
    layer2_outputs(2675) <= not((layer1_outputs(2037)) or (layer1_outputs(5629)));
    layer2_outputs(2676) <= not(layer1_outputs(2891));
    layer2_outputs(2677) <= not(layer1_outputs(4797));
    layer2_outputs(2678) <= layer1_outputs(7294);
    layer2_outputs(2679) <= layer1_outputs(2016);
    layer2_outputs(2680) <= not(layer1_outputs(9544)) or (layer1_outputs(5234));
    layer2_outputs(2681) <= not(layer1_outputs(1207));
    layer2_outputs(2682) <= not((layer1_outputs(4445)) or (layer1_outputs(8238)));
    layer2_outputs(2683) <= not(layer1_outputs(3195)) or (layer1_outputs(1487));
    layer2_outputs(2684) <= (layer1_outputs(3297)) or (layer1_outputs(5420));
    layer2_outputs(2685) <= not((layer1_outputs(5817)) xor (layer1_outputs(2237)));
    layer2_outputs(2686) <= (layer1_outputs(9431)) and not (layer1_outputs(5733));
    layer2_outputs(2687) <= not(layer1_outputs(8576));
    layer2_outputs(2688) <= not(layer1_outputs(7168));
    layer2_outputs(2689) <= not(layer1_outputs(8889));
    layer2_outputs(2690) <= not(layer1_outputs(5810));
    layer2_outputs(2691) <= layer1_outputs(2322);
    layer2_outputs(2692) <= (layer1_outputs(9633)) xor (layer1_outputs(9857));
    layer2_outputs(2693) <= (layer1_outputs(84)) and not (layer1_outputs(1858));
    layer2_outputs(2694) <= layer1_outputs(5719);
    layer2_outputs(2695) <= not(layer1_outputs(10199)) or (layer1_outputs(2427));
    layer2_outputs(2696) <= not(layer1_outputs(9219));
    layer2_outputs(2697) <= not(layer1_outputs(3382));
    layer2_outputs(2698) <= (layer1_outputs(8423)) and not (layer1_outputs(5770));
    layer2_outputs(2699) <= not((layer1_outputs(9194)) xor (layer1_outputs(7880)));
    layer2_outputs(2700) <= (layer1_outputs(2226)) xor (layer1_outputs(9412));
    layer2_outputs(2701) <= (layer1_outputs(3321)) and not (layer1_outputs(6138));
    layer2_outputs(2702) <= layer1_outputs(7605);
    layer2_outputs(2703) <= (layer1_outputs(3234)) and not (layer1_outputs(6911));
    layer2_outputs(2704) <= not((layer1_outputs(8700)) or (layer1_outputs(9955)));
    layer2_outputs(2705) <= not((layer1_outputs(3036)) and (layer1_outputs(9239)));
    layer2_outputs(2706) <= not((layer1_outputs(2168)) or (layer1_outputs(4036)));
    layer2_outputs(2707) <= not(layer1_outputs(3832));
    layer2_outputs(2708) <= not((layer1_outputs(9405)) and (layer1_outputs(381)));
    layer2_outputs(2709) <= not(layer1_outputs(3895));
    layer2_outputs(2710) <= not(layer1_outputs(8083));
    layer2_outputs(2711) <= layer1_outputs(6206);
    layer2_outputs(2712) <= not(layer1_outputs(6383));
    layer2_outputs(2713) <= not((layer1_outputs(4342)) and (layer1_outputs(2708)));
    layer2_outputs(2714) <= (layer1_outputs(5737)) or (layer1_outputs(3314));
    layer2_outputs(2715) <= layer1_outputs(9379);
    layer2_outputs(2716) <= not(layer1_outputs(4041));
    layer2_outputs(2717) <= not((layer1_outputs(4310)) xor (layer1_outputs(8891)));
    layer2_outputs(2718) <= not((layer1_outputs(2265)) xor (layer1_outputs(1673)));
    layer2_outputs(2719) <= not(layer1_outputs(9623));
    layer2_outputs(2720) <= (layer1_outputs(9423)) and not (layer1_outputs(4410));
    layer2_outputs(2721) <= not((layer1_outputs(1395)) and (layer1_outputs(9175)));
    layer2_outputs(2722) <= not((layer1_outputs(256)) or (layer1_outputs(5356)));
    layer2_outputs(2723) <= not(layer1_outputs(3597)) or (layer1_outputs(6733));
    layer2_outputs(2724) <= not((layer1_outputs(6819)) or (layer1_outputs(9655)));
    layer2_outputs(2725) <= not(layer1_outputs(3829));
    layer2_outputs(2726) <= layer1_outputs(2854);
    layer2_outputs(2727) <= not(layer1_outputs(2004));
    layer2_outputs(2728) <= (layer1_outputs(1270)) and (layer1_outputs(723));
    layer2_outputs(2729) <= not(layer1_outputs(7710)) or (layer1_outputs(9480));
    layer2_outputs(2730) <= not(layer1_outputs(9014)) or (layer1_outputs(8511));
    layer2_outputs(2731) <= not(layer1_outputs(1988));
    layer2_outputs(2732) <= (layer1_outputs(2175)) and not (layer1_outputs(9348));
    layer2_outputs(2733) <= (layer1_outputs(1700)) xor (layer1_outputs(4573));
    layer2_outputs(2734) <= (layer1_outputs(6986)) xor (layer1_outputs(1519));
    layer2_outputs(2735) <= (layer1_outputs(9044)) and not (layer1_outputs(2654));
    layer2_outputs(2736) <= not((layer1_outputs(1)) xor (layer1_outputs(7362)));
    layer2_outputs(2737) <= (layer1_outputs(257)) and not (layer1_outputs(9005));
    layer2_outputs(2738) <= layer1_outputs(5731);
    layer2_outputs(2739) <= (layer1_outputs(4776)) or (layer1_outputs(180));
    layer2_outputs(2740) <= not(layer1_outputs(3258));
    layer2_outputs(2741) <= (layer1_outputs(8264)) xor (layer1_outputs(9277));
    layer2_outputs(2742) <= layer1_outputs(7516);
    layer2_outputs(2743) <= (layer1_outputs(6517)) or (layer1_outputs(836));
    layer2_outputs(2744) <= not((layer1_outputs(5692)) and (layer1_outputs(3442)));
    layer2_outputs(2745) <= not((layer1_outputs(8563)) and (layer1_outputs(3870)));
    layer2_outputs(2746) <= not((layer1_outputs(9397)) xor (layer1_outputs(4146)));
    layer2_outputs(2747) <= not(layer1_outputs(7847));
    layer2_outputs(2748) <= not(layer1_outputs(9776));
    layer2_outputs(2749) <= layer1_outputs(8595);
    layer2_outputs(2750) <= (layer1_outputs(5173)) and (layer1_outputs(1511));
    layer2_outputs(2751) <= layer1_outputs(6510);
    layer2_outputs(2752) <= not(layer1_outputs(9165));
    layer2_outputs(2753) <= not(layer1_outputs(7614));
    layer2_outputs(2754) <= not((layer1_outputs(62)) and (layer1_outputs(6971)));
    layer2_outputs(2755) <= not(layer1_outputs(4633)) or (layer1_outputs(5540));
    layer2_outputs(2756) <= not(layer1_outputs(6963)) or (layer1_outputs(1123));
    layer2_outputs(2757) <= not(layer1_outputs(1908)) or (layer1_outputs(9403));
    layer2_outputs(2758) <= not(layer1_outputs(5988));
    layer2_outputs(2759) <= not(layer1_outputs(7297));
    layer2_outputs(2760) <= not(layer1_outputs(9635)) or (layer1_outputs(9374));
    layer2_outputs(2761) <= (layer1_outputs(8595)) and (layer1_outputs(312));
    layer2_outputs(2762) <= (layer1_outputs(7214)) and not (layer1_outputs(9438));
    layer2_outputs(2763) <= not((layer1_outputs(7789)) xor (layer1_outputs(9320)));
    layer2_outputs(2764) <= (layer1_outputs(8455)) and not (layer1_outputs(8433));
    layer2_outputs(2765) <= not((layer1_outputs(9718)) xor (layer1_outputs(1008)));
    layer2_outputs(2766) <= layer1_outputs(2078);
    layer2_outputs(2767) <= layer1_outputs(4564);
    layer2_outputs(2768) <= not(layer1_outputs(5056)) or (layer1_outputs(5609));
    layer2_outputs(2769) <= not(layer1_outputs(8445)) or (layer1_outputs(637));
    layer2_outputs(2770) <= '0';
    layer2_outputs(2771) <= layer1_outputs(3672);
    layer2_outputs(2772) <= not(layer1_outputs(10137));
    layer2_outputs(2773) <= layer1_outputs(8552);
    layer2_outputs(2774) <= (layer1_outputs(4156)) and not (layer1_outputs(8536));
    layer2_outputs(2775) <= not((layer1_outputs(5621)) and (layer1_outputs(8788)));
    layer2_outputs(2776) <= layer1_outputs(8942);
    layer2_outputs(2777) <= (layer1_outputs(6577)) and not (layer1_outputs(4603));
    layer2_outputs(2778) <= not(layer1_outputs(7369));
    layer2_outputs(2779) <= layer1_outputs(3245);
    layer2_outputs(2780) <= layer1_outputs(7692);
    layer2_outputs(2781) <= layer1_outputs(4136);
    layer2_outputs(2782) <= not((layer1_outputs(5641)) xor (layer1_outputs(5989)));
    layer2_outputs(2783) <= layer1_outputs(3800);
    layer2_outputs(2784) <= (layer1_outputs(285)) and not (layer1_outputs(8492));
    layer2_outputs(2785) <= not(layer1_outputs(2274));
    layer2_outputs(2786) <= (layer1_outputs(607)) and not (layer1_outputs(9970));
    layer2_outputs(2787) <= not((layer1_outputs(7013)) xor (layer1_outputs(1717)));
    layer2_outputs(2788) <= (layer1_outputs(841)) or (layer1_outputs(3347));
    layer2_outputs(2789) <= layer1_outputs(6543);
    layer2_outputs(2790) <= '0';
    layer2_outputs(2791) <= (layer1_outputs(1030)) and not (layer1_outputs(6703));
    layer2_outputs(2792) <= layer1_outputs(5899);
    layer2_outputs(2793) <= not((layer1_outputs(3878)) and (layer1_outputs(9946)));
    layer2_outputs(2794) <= layer1_outputs(1225);
    layer2_outputs(2795) <= not(layer1_outputs(3701));
    layer2_outputs(2796) <= not(layer1_outputs(8176));
    layer2_outputs(2797) <= (layer1_outputs(9506)) or (layer1_outputs(6848));
    layer2_outputs(2798) <= not(layer1_outputs(486));
    layer2_outputs(2799) <= layer1_outputs(1584);
    layer2_outputs(2800) <= not((layer1_outputs(7068)) xor (layer1_outputs(9482)));
    layer2_outputs(2801) <= layer1_outputs(2949);
    layer2_outputs(2802) <= layer1_outputs(8264);
    layer2_outputs(2803) <= (layer1_outputs(1460)) or (layer1_outputs(2921));
    layer2_outputs(2804) <= not(layer1_outputs(1627));
    layer2_outputs(2805) <= (layer1_outputs(5614)) and not (layer1_outputs(6439));
    layer2_outputs(2806) <= layer1_outputs(5112);
    layer2_outputs(2807) <= not(layer1_outputs(8867));
    layer2_outputs(2808) <= not(layer1_outputs(7701));
    layer2_outputs(2809) <= not(layer1_outputs(9417));
    layer2_outputs(2810) <= layer1_outputs(788);
    layer2_outputs(2811) <= (layer1_outputs(1873)) and not (layer1_outputs(969));
    layer2_outputs(2812) <= not(layer1_outputs(5534));
    layer2_outputs(2813) <= layer1_outputs(6445);
    layer2_outputs(2814) <= not((layer1_outputs(7111)) xor (layer1_outputs(813)));
    layer2_outputs(2815) <= (layer1_outputs(3853)) xor (layer1_outputs(3338));
    layer2_outputs(2816) <= not((layer1_outputs(10111)) or (layer1_outputs(2344)));
    layer2_outputs(2817) <= (layer1_outputs(1752)) and not (layer1_outputs(9826));
    layer2_outputs(2818) <= not(layer1_outputs(10102));
    layer2_outputs(2819) <= (layer1_outputs(7012)) and (layer1_outputs(511));
    layer2_outputs(2820) <= not(layer1_outputs(7960));
    layer2_outputs(2821) <= layer1_outputs(5842);
    layer2_outputs(2822) <= layer1_outputs(9619);
    layer2_outputs(2823) <= not((layer1_outputs(3086)) or (layer1_outputs(7317)));
    layer2_outputs(2824) <= (layer1_outputs(3193)) or (layer1_outputs(8259));
    layer2_outputs(2825) <= not(layer1_outputs(8136)) or (layer1_outputs(1428));
    layer2_outputs(2826) <= not(layer1_outputs(9972));
    layer2_outputs(2827) <= (layer1_outputs(7691)) or (layer1_outputs(4645));
    layer2_outputs(2828) <= not((layer1_outputs(7519)) and (layer1_outputs(1375)));
    layer2_outputs(2829) <= not(layer1_outputs(4821));
    layer2_outputs(2830) <= not((layer1_outputs(6620)) and (layer1_outputs(8320)));
    layer2_outputs(2831) <= layer1_outputs(159);
    layer2_outputs(2832) <= not(layer1_outputs(3689));
    layer2_outputs(2833) <= layer1_outputs(5886);
    layer2_outputs(2834) <= not(layer1_outputs(7605));
    layer2_outputs(2835) <= (layer1_outputs(4351)) and not (layer1_outputs(6616));
    layer2_outputs(2836) <= not(layer1_outputs(6283));
    layer2_outputs(2837) <= layer1_outputs(310);
    layer2_outputs(2838) <= layer1_outputs(5366);
    layer2_outputs(2839) <= (layer1_outputs(3976)) and not (layer1_outputs(1062));
    layer2_outputs(2840) <= not(layer1_outputs(2368));
    layer2_outputs(2841) <= not((layer1_outputs(9735)) xor (layer1_outputs(6137)));
    layer2_outputs(2842) <= not((layer1_outputs(1219)) xor (layer1_outputs(7199)));
    layer2_outputs(2843) <= (layer1_outputs(7583)) and not (layer1_outputs(7861));
    layer2_outputs(2844) <= not(layer1_outputs(5285));
    layer2_outputs(2845) <= not(layer1_outputs(3867));
    layer2_outputs(2846) <= (layer1_outputs(7957)) or (layer1_outputs(5115));
    layer2_outputs(2847) <= not(layer1_outputs(5830)) or (layer1_outputs(3254));
    layer2_outputs(2848) <= layer1_outputs(2679);
    layer2_outputs(2849) <= not(layer1_outputs(7458)) or (layer1_outputs(6273));
    layer2_outputs(2850) <= not(layer1_outputs(6479));
    layer2_outputs(2851) <= not(layer1_outputs(7956));
    layer2_outputs(2852) <= layer1_outputs(10073);
    layer2_outputs(2853) <= not(layer1_outputs(9967));
    layer2_outputs(2854) <= (layer1_outputs(7397)) and not (layer1_outputs(7773));
    layer2_outputs(2855) <= not(layer1_outputs(6981));
    layer2_outputs(2856) <= (layer1_outputs(3777)) and not (layer1_outputs(2252));
    layer2_outputs(2857) <= not((layer1_outputs(500)) and (layer1_outputs(10024)));
    layer2_outputs(2858) <= (layer1_outputs(1865)) and (layer1_outputs(7588));
    layer2_outputs(2859) <= not(layer1_outputs(7616)) or (layer1_outputs(108));
    layer2_outputs(2860) <= not((layer1_outputs(4458)) and (layer1_outputs(784)));
    layer2_outputs(2861) <= (layer1_outputs(1742)) xor (layer1_outputs(8919));
    layer2_outputs(2862) <= (layer1_outputs(7802)) and not (layer1_outputs(4032));
    layer2_outputs(2863) <= (layer1_outputs(5814)) and not (layer1_outputs(341));
    layer2_outputs(2864) <= not((layer1_outputs(1381)) or (layer1_outputs(3620)));
    layer2_outputs(2865) <= layer1_outputs(8987);
    layer2_outputs(2866) <= (layer1_outputs(3925)) and not (layer1_outputs(7492));
    layer2_outputs(2867) <= layer1_outputs(2320);
    layer2_outputs(2868) <= (layer1_outputs(5148)) or (layer1_outputs(4427));
    layer2_outputs(2869) <= layer1_outputs(6547);
    layer2_outputs(2870) <= (layer1_outputs(3945)) or (layer1_outputs(6826));
    layer2_outputs(2871) <= layer1_outputs(7556);
    layer2_outputs(2872) <= layer1_outputs(4207);
    layer2_outputs(2873) <= not((layer1_outputs(9724)) and (layer1_outputs(10104)));
    layer2_outputs(2874) <= (layer1_outputs(9656)) and not (layer1_outputs(2555));
    layer2_outputs(2875) <= not((layer1_outputs(1460)) and (layer1_outputs(6532)));
    layer2_outputs(2876) <= not((layer1_outputs(4380)) xor (layer1_outputs(2199)));
    layer2_outputs(2877) <= not((layer1_outputs(2550)) and (layer1_outputs(882)));
    layer2_outputs(2878) <= layer1_outputs(9777);
    layer2_outputs(2879) <= layer1_outputs(2469);
    layer2_outputs(2880) <= (layer1_outputs(3431)) and not (layer1_outputs(9356));
    layer2_outputs(2881) <= layer1_outputs(2331);
    layer2_outputs(2882) <= layer1_outputs(430);
    layer2_outputs(2883) <= (layer1_outputs(7792)) or (layer1_outputs(6051));
    layer2_outputs(2884) <= layer1_outputs(6639);
    layer2_outputs(2885) <= not(layer1_outputs(5235));
    layer2_outputs(2886) <= not(layer1_outputs(2815));
    layer2_outputs(2887) <= layer1_outputs(105);
    layer2_outputs(2888) <= layer1_outputs(496);
    layer2_outputs(2889) <= (layer1_outputs(5060)) and not (layer1_outputs(10017));
    layer2_outputs(2890) <= (layer1_outputs(8961)) xor (layer1_outputs(6403));
    layer2_outputs(2891) <= layer1_outputs(7694);
    layer2_outputs(2892) <= not((layer1_outputs(3111)) or (layer1_outputs(5973)));
    layer2_outputs(2893) <= (layer1_outputs(7618)) xor (layer1_outputs(10082));
    layer2_outputs(2894) <= not(layer1_outputs(7499));
    layer2_outputs(2895) <= not((layer1_outputs(7025)) xor (layer1_outputs(4368)));
    layer2_outputs(2896) <= not(layer1_outputs(9695));
    layer2_outputs(2897) <= not(layer1_outputs(6857));
    layer2_outputs(2898) <= (layer1_outputs(1640)) and not (layer1_outputs(2430));
    layer2_outputs(2899) <= not(layer1_outputs(9817));
    layer2_outputs(2900) <= (layer1_outputs(581)) and not (layer1_outputs(8015));
    layer2_outputs(2901) <= (layer1_outputs(9406)) and (layer1_outputs(7758));
    layer2_outputs(2902) <= not((layer1_outputs(7354)) or (layer1_outputs(7829)));
    layer2_outputs(2903) <= not(layer1_outputs(3513));
    layer2_outputs(2904) <= layer1_outputs(514);
    layer2_outputs(2905) <= not((layer1_outputs(2576)) and (layer1_outputs(5152)));
    layer2_outputs(2906) <= layer1_outputs(5603);
    layer2_outputs(2907) <= (layer1_outputs(4097)) and not (layer1_outputs(3167));
    layer2_outputs(2908) <= not((layer1_outputs(2618)) xor (layer1_outputs(8285)));
    layer2_outputs(2909) <= (layer1_outputs(6367)) and not (layer1_outputs(8042));
    layer2_outputs(2910) <= not(layer1_outputs(768));
    layer2_outputs(2911) <= '0';
    layer2_outputs(2912) <= layer1_outputs(9540);
    layer2_outputs(2913) <= (layer1_outputs(7958)) or (layer1_outputs(10121));
    layer2_outputs(2914) <= (layer1_outputs(3788)) and not (layer1_outputs(8315));
    layer2_outputs(2915) <= (layer1_outputs(2932)) or (layer1_outputs(6659));
    layer2_outputs(2916) <= layer1_outputs(2712);
    layer2_outputs(2917) <= (layer1_outputs(6618)) and not (layer1_outputs(8078));
    layer2_outputs(2918) <= not(layer1_outputs(5982)) or (layer1_outputs(584));
    layer2_outputs(2919) <= (layer1_outputs(3640)) and not (layer1_outputs(2557));
    layer2_outputs(2920) <= not(layer1_outputs(9435));
    layer2_outputs(2921) <= not(layer1_outputs(6396));
    layer2_outputs(2922) <= not(layer1_outputs(5704));
    layer2_outputs(2923) <= not(layer1_outputs(1753));
    layer2_outputs(2924) <= not(layer1_outputs(8492));
    layer2_outputs(2925) <= not(layer1_outputs(6066)) or (layer1_outputs(7681));
    layer2_outputs(2926) <= not((layer1_outputs(4630)) or (layer1_outputs(1957)));
    layer2_outputs(2927) <= layer1_outputs(2975);
    layer2_outputs(2928) <= layer1_outputs(10140);
    layer2_outputs(2929) <= (layer1_outputs(846)) xor (layer1_outputs(9736));
    layer2_outputs(2930) <= (layer1_outputs(9696)) xor (layer1_outputs(3926));
    layer2_outputs(2931) <= not(layer1_outputs(6706)) or (layer1_outputs(1845));
    layer2_outputs(2932) <= layer1_outputs(5260);
    layer2_outputs(2933) <= not((layer1_outputs(7106)) or (layer1_outputs(2082)));
    layer2_outputs(2934) <= not(layer1_outputs(3155)) or (layer1_outputs(917));
    layer2_outputs(2935) <= not((layer1_outputs(6511)) xor (layer1_outputs(7320)));
    layer2_outputs(2936) <= (layer1_outputs(3413)) and (layer1_outputs(3179));
    layer2_outputs(2937) <= (layer1_outputs(9855)) and (layer1_outputs(2002));
    layer2_outputs(2938) <= not(layer1_outputs(6194));
    layer2_outputs(2939) <= not(layer1_outputs(5583));
    layer2_outputs(2940) <= not(layer1_outputs(9746));
    layer2_outputs(2941) <= (layer1_outputs(7612)) xor (layer1_outputs(5584));
    layer2_outputs(2942) <= (layer1_outputs(10054)) and not (layer1_outputs(6043));
    layer2_outputs(2943) <= (layer1_outputs(233)) and not (layer1_outputs(678));
    layer2_outputs(2944) <= layer1_outputs(3503);
    layer2_outputs(2945) <= not(layer1_outputs(7256));
    layer2_outputs(2946) <= not(layer1_outputs(7189)) or (layer1_outputs(8061));
    layer2_outputs(2947) <= not(layer1_outputs(2916));
    layer2_outputs(2948) <= not((layer1_outputs(4691)) xor (layer1_outputs(455)));
    layer2_outputs(2949) <= (layer1_outputs(6544)) and (layer1_outputs(5656));
    layer2_outputs(2950) <= (layer1_outputs(2935)) xor (layer1_outputs(143));
    layer2_outputs(2951) <= (layer1_outputs(5846)) and not (layer1_outputs(5843));
    layer2_outputs(2952) <= not((layer1_outputs(7445)) xor (layer1_outputs(7505)));
    layer2_outputs(2953) <= not(layer1_outputs(386));
    layer2_outputs(2954) <= not(layer1_outputs(7211)) or (layer1_outputs(9322));
    layer2_outputs(2955) <= (layer1_outputs(3621)) and (layer1_outputs(8596));
    layer2_outputs(2956) <= (layer1_outputs(698)) and not (layer1_outputs(3349));
    layer2_outputs(2957) <= not(layer1_outputs(301));
    layer2_outputs(2958) <= not(layer1_outputs(6730));
    layer2_outputs(2959) <= not((layer1_outputs(8294)) xor (layer1_outputs(2903)));
    layer2_outputs(2960) <= not(layer1_outputs(6995)) or (layer1_outputs(386));
    layer2_outputs(2961) <= '0';
    layer2_outputs(2962) <= layer1_outputs(925);
    layer2_outputs(2963) <= layer1_outputs(2433);
    layer2_outputs(2964) <= not((layer1_outputs(4078)) xor (layer1_outputs(2686)));
    layer2_outputs(2965) <= (layer1_outputs(2348)) and not (layer1_outputs(7994));
    layer2_outputs(2966) <= not(layer1_outputs(7799));
    layer2_outputs(2967) <= (layer1_outputs(1330)) and not (layer1_outputs(1977));
    layer2_outputs(2968) <= not((layer1_outputs(5923)) or (layer1_outputs(9741)));
    layer2_outputs(2969) <= (layer1_outputs(7904)) or (layer1_outputs(4585));
    layer2_outputs(2970) <= layer1_outputs(6295);
    layer2_outputs(2971) <= not(layer1_outputs(3276)) or (layer1_outputs(2198));
    layer2_outputs(2972) <= (layer1_outputs(5953)) and not (layer1_outputs(4720));
    layer2_outputs(2973) <= not(layer1_outputs(2098));
    layer2_outputs(2974) <= not(layer1_outputs(6401)) or (layer1_outputs(2896));
    layer2_outputs(2975) <= not(layer1_outputs(2050));
    layer2_outputs(2976) <= layer1_outputs(465);
    layer2_outputs(2977) <= not(layer1_outputs(7138));
    layer2_outputs(2978) <= layer1_outputs(6167);
    layer2_outputs(2979) <= not(layer1_outputs(8555));
    layer2_outputs(2980) <= layer1_outputs(1370);
    layer2_outputs(2981) <= layer1_outputs(4859);
    layer2_outputs(2982) <= not(layer1_outputs(7028));
    layer2_outputs(2983) <= not((layer1_outputs(2111)) and (layer1_outputs(8385)));
    layer2_outputs(2984) <= not(layer1_outputs(9284));
    layer2_outputs(2985) <= (layer1_outputs(10204)) or (layer1_outputs(4110));
    layer2_outputs(2986) <= (layer1_outputs(9761)) or (layer1_outputs(7720));
    layer2_outputs(2987) <= layer1_outputs(8968);
    layer2_outputs(2988) <= not(layer1_outputs(3446)) or (layer1_outputs(856));
    layer2_outputs(2989) <= layer1_outputs(101);
    layer2_outputs(2990) <= not(layer1_outputs(8882)) or (layer1_outputs(9583));
    layer2_outputs(2991) <= layer1_outputs(2706);
    layer2_outputs(2992) <= not(layer1_outputs(7292));
    layer2_outputs(2993) <= not((layer1_outputs(4494)) and (layer1_outputs(6437)));
    layer2_outputs(2994) <= not((layer1_outputs(1726)) xor (layer1_outputs(3192)));
    layer2_outputs(2995) <= not(layer1_outputs(4383));
    layer2_outputs(2996) <= layer1_outputs(6865);
    layer2_outputs(2997) <= layer1_outputs(2020);
    layer2_outputs(2998) <= not((layer1_outputs(2353)) and (layer1_outputs(6637)));
    layer2_outputs(2999) <= layer1_outputs(9800);
    layer2_outputs(3000) <= not(layer1_outputs(1500)) or (layer1_outputs(10103));
    layer2_outputs(3001) <= (layer1_outputs(7315)) xor (layer1_outputs(8018));
    layer2_outputs(3002) <= (layer1_outputs(6947)) xor (layer1_outputs(10054));
    layer2_outputs(3003) <= (layer1_outputs(6850)) and (layer1_outputs(8854));
    layer2_outputs(3004) <= (layer1_outputs(4200)) xor (layer1_outputs(9906));
    layer2_outputs(3005) <= not(layer1_outputs(2454)) or (layer1_outputs(1601));
    layer2_outputs(3006) <= not(layer1_outputs(8890)) or (layer1_outputs(1207));
    layer2_outputs(3007) <= not((layer1_outputs(1724)) xor (layer1_outputs(7985)));
    layer2_outputs(3008) <= (layer1_outputs(1070)) or (layer1_outputs(5960));
    layer2_outputs(3009) <= not(layer1_outputs(344));
    layer2_outputs(3010) <= layer1_outputs(2135);
    layer2_outputs(3011) <= not(layer1_outputs(645));
    layer2_outputs(3012) <= layer1_outputs(9732);
    layer2_outputs(3013) <= not((layer1_outputs(9677)) xor (layer1_outputs(7545)));
    layer2_outputs(3014) <= (layer1_outputs(6938)) and (layer1_outputs(5353));
    layer2_outputs(3015) <= layer1_outputs(8833);
    layer2_outputs(3016) <= layer1_outputs(3970);
    layer2_outputs(3017) <= not(layer1_outputs(6845));
    layer2_outputs(3018) <= not((layer1_outputs(3200)) xor (layer1_outputs(3837)));
    layer2_outputs(3019) <= not(layer1_outputs(4852));
    layer2_outputs(3020) <= not((layer1_outputs(6119)) and (layer1_outputs(6494)));
    layer2_outputs(3021) <= not((layer1_outputs(9944)) xor (layer1_outputs(9649)));
    layer2_outputs(3022) <= (layer1_outputs(6106)) and not (layer1_outputs(760));
    layer2_outputs(3023) <= (layer1_outputs(3363)) or (layer1_outputs(2616));
    layer2_outputs(3024) <= not(layer1_outputs(10103)) or (layer1_outputs(8487));
    layer2_outputs(3025) <= not((layer1_outputs(4084)) xor (layer1_outputs(3820)));
    layer2_outputs(3026) <= not(layer1_outputs(8189));
    layer2_outputs(3027) <= not(layer1_outputs(6228));
    layer2_outputs(3028) <= (layer1_outputs(9478)) or (layer1_outputs(8203));
    layer2_outputs(3029) <= (layer1_outputs(4857)) and not (layer1_outputs(747));
    layer2_outputs(3030) <= not(layer1_outputs(5680));
    layer2_outputs(3031) <= not(layer1_outputs(1852));
    layer2_outputs(3032) <= layer1_outputs(1995);
    layer2_outputs(3033) <= not(layer1_outputs(7883));
    layer2_outputs(3034) <= not(layer1_outputs(4387));
    layer2_outputs(3035) <= layer1_outputs(313);
    layer2_outputs(3036) <= (layer1_outputs(1891)) and not (layer1_outputs(6351));
    layer2_outputs(3037) <= not((layer1_outputs(1664)) xor (layer1_outputs(5713)));
    layer2_outputs(3038) <= not(layer1_outputs(541)) or (layer1_outputs(7283));
    layer2_outputs(3039) <= (layer1_outputs(4668)) and (layer1_outputs(5952));
    layer2_outputs(3040) <= (layer1_outputs(10172)) and (layer1_outputs(6198));
    layer2_outputs(3041) <= not(layer1_outputs(7653)) or (layer1_outputs(3679));
    layer2_outputs(3042) <= not(layer1_outputs(7428));
    layer2_outputs(3043) <= layer1_outputs(217);
    layer2_outputs(3044) <= not((layer1_outputs(7845)) or (layer1_outputs(1644)));
    layer2_outputs(3045) <= not(layer1_outputs(5881));
    layer2_outputs(3046) <= layer1_outputs(3998);
    layer2_outputs(3047) <= not(layer1_outputs(2293));
    layer2_outputs(3048) <= not((layer1_outputs(2620)) and (layer1_outputs(6263)));
    layer2_outputs(3049) <= not((layer1_outputs(8321)) xor (layer1_outputs(9796)));
    layer2_outputs(3050) <= not(layer1_outputs(8980));
    layer2_outputs(3051) <= (layer1_outputs(3018)) and not (layer1_outputs(4373));
    layer2_outputs(3052) <= not(layer1_outputs(8160));
    layer2_outputs(3053) <= not(layer1_outputs(4040));
    layer2_outputs(3054) <= (layer1_outputs(811)) xor (layer1_outputs(2434));
    layer2_outputs(3055) <= layer1_outputs(5711);
    layer2_outputs(3056) <= not(layer1_outputs(2455));
    layer2_outputs(3057) <= not(layer1_outputs(421));
    layer2_outputs(3058) <= layer1_outputs(9247);
    layer2_outputs(3059) <= not(layer1_outputs(7114));
    layer2_outputs(3060) <= not((layer1_outputs(2141)) and (layer1_outputs(3657)));
    layer2_outputs(3061) <= not(layer1_outputs(3201));
    layer2_outputs(3062) <= not(layer1_outputs(169)) or (layer1_outputs(9901));
    layer2_outputs(3063) <= not(layer1_outputs(9310));
    layer2_outputs(3064) <= not(layer1_outputs(2601)) or (layer1_outputs(4721));
    layer2_outputs(3065) <= (layer1_outputs(7875)) and not (layer1_outputs(9144));
    layer2_outputs(3066) <= not((layer1_outputs(1459)) and (layer1_outputs(9300)));
    layer2_outputs(3067) <= (layer1_outputs(2869)) xor (layer1_outputs(2443));
    layer2_outputs(3068) <= not(layer1_outputs(7011));
    layer2_outputs(3069) <= not(layer1_outputs(6054));
    layer2_outputs(3070) <= not(layer1_outputs(5943));
    layer2_outputs(3071) <= not(layer1_outputs(3165));
    layer2_outputs(3072) <= layer1_outputs(4536);
    layer2_outputs(3073) <= not(layer1_outputs(6392));
    layer2_outputs(3074) <= (layer1_outputs(6565)) xor (layer1_outputs(2201));
    layer2_outputs(3075) <= not(layer1_outputs(4198));
    layer2_outputs(3076) <= layer1_outputs(4614);
    layer2_outputs(3077) <= not((layer1_outputs(2962)) or (layer1_outputs(10101)));
    layer2_outputs(3078) <= (layer1_outputs(9627)) xor (layer1_outputs(2230));
    layer2_outputs(3079) <= not((layer1_outputs(4253)) and (layer1_outputs(7375)));
    layer2_outputs(3080) <= not(layer1_outputs(8008));
    layer2_outputs(3081) <= not(layer1_outputs(221));
    layer2_outputs(3082) <= not((layer1_outputs(9603)) xor (layer1_outputs(9418)));
    layer2_outputs(3083) <= not(layer1_outputs(5977)) or (layer1_outputs(9565));
    layer2_outputs(3084) <= not((layer1_outputs(4498)) and (layer1_outputs(4900)));
    layer2_outputs(3085) <= (layer1_outputs(2997)) xor (layer1_outputs(2527));
    layer2_outputs(3086) <= (layer1_outputs(6531)) xor (layer1_outputs(574));
    layer2_outputs(3087) <= layer1_outputs(4751);
    layer2_outputs(3088) <= '0';
    layer2_outputs(3089) <= not((layer1_outputs(4383)) or (layer1_outputs(9452)));
    layer2_outputs(3090) <= not((layer1_outputs(10015)) and (layer1_outputs(8333)));
    layer2_outputs(3091) <= not((layer1_outputs(941)) xor (layer1_outputs(8795)));
    layer2_outputs(3092) <= not((layer1_outputs(7595)) and (layer1_outputs(1636)));
    layer2_outputs(3093) <= not(layer1_outputs(6648)) or (layer1_outputs(3198));
    layer2_outputs(3094) <= (layer1_outputs(2306)) and (layer1_outputs(4102));
    layer2_outputs(3095) <= (layer1_outputs(9299)) and not (layer1_outputs(9528));
    layer2_outputs(3096) <= (layer1_outputs(9432)) and (layer1_outputs(1762));
    layer2_outputs(3097) <= not(layer1_outputs(8183)) or (layer1_outputs(3487));
    layer2_outputs(3098) <= layer1_outputs(6688);
    layer2_outputs(3099) <= not((layer1_outputs(3093)) or (layer1_outputs(9922)));
    layer2_outputs(3100) <= layer1_outputs(962);
    layer2_outputs(3101) <= not(layer1_outputs(7830));
    layer2_outputs(3102) <= layer1_outputs(3705);
    layer2_outputs(3103) <= not(layer1_outputs(8118)) or (layer1_outputs(715));
    layer2_outputs(3104) <= not((layer1_outputs(6366)) or (layer1_outputs(7153)));
    layer2_outputs(3105) <= layer1_outputs(2895);
    layer2_outputs(3106) <= layer1_outputs(10055);
    layer2_outputs(3107) <= not(layer1_outputs(3826));
    layer2_outputs(3108) <= (layer1_outputs(636)) and not (layer1_outputs(9336));
    layer2_outputs(3109) <= layer1_outputs(8269);
    layer2_outputs(3110) <= layer1_outputs(1658);
    layer2_outputs(3111) <= not(layer1_outputs(9557));
    layer2_outputs(3112) <= not(layer1_outputs(1981));
    layer2_outputs(3113) <= not(layer1_outputs(4348));
    layer2_outputs(3114) <= not(layer1_outputs(2254));
    layer2_outputs(3115) <= not(layer1_outputs(3963));
    layer2_outputs(3116) <= layer1_outputs(6528);
    layer2_outputs(3117) <= not(layer1_outputs(2894)) or (layer1_outputs(9498));
    layer2_outputs(3118) <= not(layer1_outputs(609));
    layer2_outputs(3119) <= not(layer1_outputs(7676));
    layer2_outputs(3120) <= not(layer1_outputs(3417)) or (layer1_outputs(9346));
    layer2_outputs(3121) <= not((layer1_outputs(320)) and (layer1_outputs(2318)));
    layer2_outputs(3122) <= not(layer1_outputs(358)) or (layer1_outputs(7116));
    layer2_outputs(3123) <= not(layer1_outputs(6890));
    layer2_outputs(3124) <= not(layer1_outputs(1837));
    layer2_outputs(3125) <= layer1_outputs(7203);
    layer2_outputs(3126) <= layer1_outputs(1357);
    layer2_outputs(3127) <= not(layer1_outputs(4461)) or (layer1_outputs(6929));
    layer2_outputs(3128) <= layer1_outputs(5105);
    layer2_outputs(3129) <= not((layer1_outputs(7821)) xor (layer1_outputs(7582)));
    layer2_outputs(3130) <= not(layer1_outputs(2541));
    layer2_outputs(3131) <= not((layer1_outputs(7347)) and (layer1_outputs(6714)));
    layer2_outputs(3132) <= not(layer1_outputs(8738));
    layer2_outputs(3133) <= not(layer1_outputs(5101));
    layer2_outputs(3134) <= not(layer1_outputs(1416));
    layer2_outputs(3135) <= not(layer1_outputs(8666));
    layer2_outputs(3136) <= (layer1_outputs(9019)) xor (layer1_outputs(1481));
    layer2_outputs(3137) <= not(layer1_outputs(7214));
    layer2_outputs(3138) <= layer1_outputs(6346);
    layer2_outputs(3139) <= layer1_outputs(3994);
    layer2_outputs(3140) <= (layer1_outputs(702)) and not (layer1_outputs(517));
    layer2_outputs(3141) <= not((layer1_outputs(2881)) or (layer1_outputs(2171)));
    layer2_outputs(3142) <= (layer1_outputs(6785)) and not (layer1_outputs(3089));
    layer2_outputs(3143) <= not(layer1_outputs(8735));
    layer2_outputs(3144) <= not(layer1_outputs(9045));
    layer2_outputs(3145) <= not(layer1_outputs(8906));
    layer2_outputs(3146) <= not(layer1_outputs(5315));
    layer2_outputs(3147) <= not((layer1_outputs(1952)) xor (layer1_outputs(3681)));
    layer2_outputs(3148) <= not(layer1_outputs(7929));
    layer2_outputs(3149) <= (layer1_outputs(2110)) and not (layer1_outputs(6953));
    layer2_outputs(3150) <= not(layer1_outputs(3315)) or (layer1_outputs(2629));
    layer2_outputs(3151) <= layer1_outputs(8639);
    layer2_outputs(3152) <= layer1_outputs(6504);
    layer2_outputs(3153) <= not((layer1_outputs(4291)) or (layer1_outputs(2224)));
    layer2_outputs(3154) <= layer1_outputs(612);
    layer2_outputs(3155) <= not((layer1_outputs(5699)) and (layer1_outputs(5139)));
    layer2_outputs(3156) <= not(layer1_outputs(5083));
    layer2_outputs(3157) <= (layer1_outputs(1644)) xor (layer1_outputs(8241));
    layer2_outputs(3158) <= layer1_outputs(8489);
    layer2_outputs(3159) <= (layer1_outputs(2166)) xor (layer1_outputs(4192));
    layer2_outputs(3160) <= not(layer1_outputs(1985));
    layer2_outputs(3161) <= layer1_outputs(4814);
    layer2_outputs(3162) <= not(layer1_outputs(3063));
    layer2_outputs(3163) <= not(layer1_outputs(7049));
    layer2_outputs(3164) <= not(layer1_outputs(5170)) or (layer1_outputs(2579));
    layer2_outputs(3165) <= layer1_outputs(9034);
    layer2_outputs(3166) <= not(layer1_outputs(1985));
    layer2_outputs(3167) <= not(layer1_outputs(6529)) or (layer1_outputs(7935));
    layer2_outputs(3168) <= not(layer1_outputs(7272));
    layer2_outputs(3169) <= not(layer1_outputs(2303)) or (layer1_outputs(8953));
    layer2_outputs(3170) <= not(layer1_outputs(5973)) or (layer1_outputs(7289));
    layer2_outputs(3171) <= layer1_outputs(2211);
    layer2_outputs(3172) <= not((layer1_outputs(8125)) or (layer1_outputs(7077)));
    layer2_outputs(3173) <= not(layer1_outputs(8395));
    layer2_outputs(3174) <= not(layer1_outputs(2247));
    layer2_outputs(3175) <= not(layer1_outputs(213));
    layer2_outputs(3176) <= not(layer1_outputs(6744));
    layer2_outputs(3177) <= not(layer1_outputs(9772)) or (layer1_outputs(9379));
    layer2_outputs(3178) <= not((layer1_outputs(9298)) and (layer1_outputs(3903)));
    layer2_outputs(3179) <= not(layer1_outputs(1721));
    layer2_outputs(3180) <= not(layer1_outputs(5055));
    layer2_outputs(3181) <= not(layer1_outputs(1968)) or (layer1_outputs(10217));
    layer2_outputs(3182) <= not(layer1_outputs(8456));
    layer2_outputs(3183) <= layer1_outputs(2972);
    layer2_outputs(3184) <= layer1_outputs(5947);
    layer2_outputs(3185) <= layer1_outputs(8601);
    layer2_outputs(3186) <= not(layer1_outputs(3339));
    layer2_outputs(3187) <= layer1_outputs(6337);
    layer2_outputs(3188) <= not(layer1_outputs(549));
    layer2_outputs(3189) <= (layer1_outputs(4470)) or (layer1_outputs(6573));
    layer2_outputs(3190) <= not(layer1_outputs(5611));
    layer2_outputs(3191) <= (layer1_outputs(1749)) xor (layer1_outputs(4343));
    layer2_outputs(3192) <= not(layer1_outputs(7275)) or (layer1_outputs(1765));
    layer2_outputs(3193) <= (layer1_outputs(5958)) and not (layer1_outputs(2293));
    layer2_outputs(3194) <= not((layer1_outputs(7796)) and (layer1_outputs(2524)));
    layer2_outputs(3195) <= not(layer1_outputs(7378));
    layer2_outputs(3196) <= not(layer1_outputs(1928));
    layer2_outputs(3197) <= not(layer1_outputs(2461)) or (layer1_outputs(8760));
    layer2_outputs(3198) <= not(layer1_outputs(3028));
    layer2_outputs(3199) <= layer1_outputs(6530);
    layer2_outputs(3200) <= not(layer1_outputs(9809)) or (layer1_outputs(8195));
    layer2_outputs(3201) <= (layer1_outputs(2617)) xor (layer1_outputs(113));
    layer2_outputs(3202) <= (layer1_outputs(9094)) and (layer1_outputs(9081));
    layer2_outputs(3203) <= (layer1_outputs(7626)) and not (layer1_outputs(153));
    layer2_outputs(3204) <= (layer1_outputs(9041)) and (layer1_outputs(3972));
    layer2_outputs(3205) <= not((layer1_outputs(498)) and (layer1_outputs(6485)));
    layer2_outputs(3206) <= (layer1_outputs(5031)) xor (layer1_outputs(1810));
    layer2_outputs(3207) <= not(layer1_outputs(9663));
    layer2_outputs(3208) <= (layer1_outputs(5294)) and not (layer1_outputs(6664));
    layer2_outputs(3209) <= layer1_outputs(5998);
    layer2_outputs(3210) <= not(layer1_outputs(9816));
    layer2_outputs(3211) <= layer1_outputs(2596);
    layer2_outputs(3212) <= (layer1_outputs(5757)) and (layer1_outputs(2053));
    layer2_outputs(3213) <= (layer1_outputs(2948)) xor (layer1_outputs(4491));
    layer2_outputs(3214) <= layer1_outputs(7610);
    layer2_outputs(3215) <= not(layer1_outputs(10040));
    layer2_outputs(3216) <= not((layer1_outputs(508)) and (layer1_outputs(5542)));
    layer2_outputs(3217) <= not((layer1_outputs(6512)) and (layer1_outputs(6587)));
    layer2_outputs(3218) <= not(layer1_outputs(9636));
    layer2_outputs(3219) <= layer1_outputs(7623);
    layer2_outputs(3220) <= (layer1_outputs(5374)) and not (layer1_outputs(8566));
    layer2_outputs(3221) <= not((layer1_outputs(1982)) xor (layer1_outputs(6358)));
    layer2_outputs(3222) <= (layer1_outputs(6540)) and (layer1_outputs(4155));
    layer2_outputs(3223) <= layer1_outputs(9439);
    layer2_outputs(3224) <= (layer1_outputs(6971)) and not (layer1_outputs(4482));
    layer2_outputs(3225) <= (layer1_outputs(5049)) xor (layer1_outputs(4903));
    layer2_outputs(3226) <= not((layer1_outputs(2904)) or (layer1_outputs(4101)));
    layer2_outputs(3227) <= (layer1_outputs(9264)) or (layer1_outputs(7453));
    layer2_outputs(3228) <= layer1_outputs(4564);
    layer2_outputs(3229) <= not(layer1_outputs(9695));
    layer2_outputs(3230) <= (layer1_outputs(3039)) or (layer1_outputs(823));
    layer2_outputs(3231) <= not(layer1_outputs(2181));
    layer2_outputs(3232) <= (layer1_outputs(6186)) and not (layer1_outputs(9639));
    layer2_outputs(3233) <= layer1_outputs(9223);
    layer2_outputs(3234) <= (layer1_outputs(1648)) and (layer1_outputs(6802));
    layer2_outputs(3235) <= layer1_outputs(2890);
    layer2_outputs(3236) <= not((layer1_outputs(3509)) and (layer1_outputs(5955)));
    layer2_outputs(3237) <= (layer1_outputs(6088)) and not (layer1_outputs(5980));
    layer2_outputs(3238) <= not(layer1_outputs(5532)) or (layer1_outputs(3298));
    layer2_outputs(3239) <= not(layer1_outputs(3397));
    layer2_outputs(3240) <= (layer1_outputs(7675)) and not (layer1_outputs(4693));
    layer2_outputs(3241) <= layer1_outputs(7725);
    layer2_outputs(3242) <= not((layer1_outputs(10049)) and (layer1_outputs(9769)));
    layer2_outputs(3243) <= not((layer1_outputs(9748)) xor (layer1_outputs(8436)));
    layer2_outputs(3244) <= not(layer1_outputs(7822));
    layer2_outputs(3245) <= not(layer1_outputs(6713));
    layer2_outputs(3246) <= not(layer1_outputs(3849));
    layer2_outputs(3247) <= (layer1_outputs(1400)) and (layer1_outputs(9205));
    layer2_outputs(3248) <= layer1_outputs(1261);
    layer2_outputs(3249) <= (layer1_outputs(2672)) or (layer1_outputs(7362));
    layer2_outputs(3250) <= layer1_outputs(1621);
    layer2_outputs(3251) <= not(layer1_outputs(5156)) or (layer1_outputs(9236));
    layer2_outputs(3252) <= not(layer1_outputs(149));
    layer2_outputs(3253) <= not(layer1_outputs(1019));
    layer2_outputs(3254) <= layer1_outputs(1545);
    layer2_outputs(3255) <= (layer1_outputs(10085)) and not (layer1_outputs(10023));
    layer2_outputs(3256) <= (layer1_outputs(3932)) and (layer1_outputs(92));
    layer2_outputs(3257) <= not(layer1_outputs(5730));
    layer2_outputs(3258) <= layer1_outputs(6871);
    layer2_outputs(3259) <= not(layer1_outputs(3548)) or (layer1_outputs(2753));
    layer2_outputs(3260) <= not(layer1_outputs(4323));
    layer2_outputs(3261) <= layer1_outputs(3574);
    layer2_outputs(3262) <= '1';
    layer2_outputs(3263) <= (layer1_outputs(3049)) or (layer1_outputs(8675));
    layer2_outputs(3264) <= (layer1_outputs(4744)) and not (layer1_outputs(142));
    layer2_outputs(3265) <= (layer1_outputs(8155)) and not (layer1_outputs(817));
    layer2_outputs(3266) <= (layer1_outputs(62)) xor (layer1_outputs(7464));
    layer2_outputs(3267) <= not((layer1_outputs(9813)) or (layer1_outputs(2641)));
    layer2_outputs(3268) <= not((layer1_outputs(993)) and (layer1_outputs(6766)));
    layer2_outputs(3269) <= not((layer1_outputs(1382)) xor (layer1_outputs(5062)));
    layer2_outputs(3270) <= not(layer1_outputs(1080));
    layer2_outputs(3271) <= not(layer1_outputs(6204));
    layer2_outputs(3272) <= (layer1_outputs(8173)) xor (layer1_outputs(4568));
    layer2_outputs(3273) <= (layer1_outputs(1149)) and (layer1_outputs(597));
    layer2_outputs(3274) <= layer1_outputs(3458);
    layer2_outputs(3275) <= not(layer1_outputs(3626));
    layer2_outputs(3276) <= layer1_outputs(2242);
    layer2_outputs(3277) <= not(layer1_outputs(10031)) or (layer1_outputs(7215));
    layer2_outputs(3278) <= layer1_outputs(6982);
    layer2_outputs(3279) <= '0';
    layer2_outputs(3280) <= layer1_outputs(1469);
    layer2_outputs(3281) <= not((layer1_outputs(6738)) or (layer1_outputs(2289)));
    layer2_outputs(3282) <= not(layer1_outputs(4322));
    layer2_outputs(3283) <= layer1_outputs(3749);
    layer2_outputs(3284) <= not(layer1_outputs(2070));
    layer2_outputs(3285) <= not(layer1_outputs(8888));
    layer2_outputs(3286) <= (layer1_outputs(7704)) or (layer1_outputs(290));
    layer2_outputs(3287) <= not(layer1_outputs(1057)) or (layer1_outputs(2766));
    layer2_outputs(3288) <= not(layer1_outputs(3441)) or (layer1_outputs(2139));
    layer2_outputs(3289) <= not((layer1_outputs(2281)) or (layer1_outputs(9214)));
    layer2_outputs(3290) <= not((layer1_outputs(9135)) xor (layer1_outputs(9144)));
    layer2_outputs(3291) <= not(layer1_outputs(1295)) or (layer1_outputs(427));
    layer2_outputs(3292) <= (layer1_outputs(8465)) and not (layer1_outputs(958));
    layer2_outputs(3293) <= (layer1_outputs(9105)) xor (layer1_outputs(9521));
    layer2_outputs(3294) <= not(layer1_outputs(9225));
    layer2_outputs(3295) <= (layer1_outputs(2613)) and (layer1_outputs(9653));
    layer2_outputs(3296) <= (layer1_outputs(6232)) and (layer1_outputs(7993));
    layer2_outputs(3297) <= not((layer1_outputs(7996)) xor (layer1_outputs(419)));
    layer2_outputs(3298) <= '1';
    layer2_outputs(3299) <= layer1_outputs(4727);
    layer2_outputs(3300) <= not(layer1_outputs(6682));
    layer2_outputs(3301) <= not(layer1_outputs(8291));
    layer2_outputs(3302) <= layer1_outputs(9147);
    layer2_outputs(3303) <= not((layer1_outputs(3570)) xor (layer1_outputs(4598)));
    layer2_outputs(3304) <= not(layer1_outputs(8292));
    layer2_outputs(3305) <= not((layer1_outputs(6431)) and (layer1_outputs(3721)));
    layer2_outputs(3306) <= (layer1_outputs(8473)) or (layer1_outputs(6781));
    layer2_outputs(3307) <= layer1_outputs(3205);
    layer2_outputs(3308) <= (layer1_outputs(8096)) and (layer1_outputs(4566));
    layer2_outputs(3309) <= not((layer1_outputs(6527)) and (layer1_outputs(8822)));
    layer2_outputs(3310) <= not(layer1_outputs(8602)) or (layer1_outputs(6169));
    layer2_outputs(3311) <= not((layer1_outputs(10232)) and (layer1_outputs(9534)));
    layer2_outputs(3312) <= not((layer1_outputs(4682)) or (layer1_outputs(219)));
    layer2_outputs(3313) <= not(layer1_outputs(4025));
    layer2_outputs(3314) <= not(layer1_outputs(6830));
    layer2_outputs(3315) <= layer1_outputs(6311);
    layer2_outputs(3316) <= not(layer1_outputs(10013));
    layer2_outputs(3317) <= not(layer1_outputs(994));
    layer2_outputs(3318) <= not(layer1_outputs(6737));
    layer2_outputs(3319) <= not(layer1_outputs(4177));
    layer2_outputs(3320) <= not((layer1_outputs(9284)) and (layer1_outputs(845)));
    layer2_outputs(3321) <= not(layer1_outputs(1242)) or (layer1_outputs(7014));
    layer2_outputs(3322) <= (layer1_outputs(2389)) and (layer1_outputs(489));
    layer2_outputs(3323) <= not(layer1_outputs(9046));
    layer2_outputs(3324) <= (layer1_outputs(4589)) and not (layer1_outputs(3430));
    layer2_outputs(3325) <= not(layer1_outputs(3879));
    layer2_outputs(3326) <= (layer1_outputs(8545)) and (layer1_outputs(2828));
    layer2_outputs(3327) <= (layer1_outputs(3439)) and not (layer1_outputs(9118));
    layer2_outputs(3328) <= layer1_outputs(7542);
    layer2_outputs(3329) <= not((layer1_outputs(7977)) xor (layer1_outputs(6356)));
    layer2_outputs(3330) <= (layer1_outputs(9514)) and not (layer1_outputs(1142));
    layer2_outputs(3331) <= (layer1_outputs(1959)) or (layer1_outputs(4365));
    layer2_outputs(3332) <= not((layer1_outputs(9336)) xor (layer1_outputs(7627)));
    layer2_outputs(3333) <= (layer1_outputs(9597)) and not (layer1_outputs(9268));
    layer2_outputs(3334) <= not((layer1_outputs(6075)) xor (layer1_outputs(5359)));
    layer2_outputs(3335) <= not(layer1_outputs(10122));
    layer2_outputs(3336) <= layer1_outputs(5421);
    layer2_outputs(3337) <= (layer1_outputs(3902)) and not (layer1_outputs(3412));
    layer2_outputs(3338) <= not(layer1_outputs(9688));
    layer2_outputs(3339) <= not(layer1_outputs(4629));
    layer2_outputs(3340) <= layer1_outputs(68);
    layer2_outputs(3341) <= layer1_outputs(9821);
    layer2_outputs(3342) <= not(layer1_outputs(3027)) or (layer1_outputs(7969));
    layer2_outputs(3343) <= not((layer1_outputs(9496)) or (layer1_outputs(1827)));
    layer2_outputs(3344) <= (layer1_outputs(4766)) xor (layer1_outputs(6651));
    layer2_outputs(3345) <= layer1_outputs(7842);
    layer2_outputs(3346) <= not(layer1_outputs(7391)) or (layer1_outputs(6021));
    layer2_outputs(3347) <= not((layer1_outputs(1971)) or (layer1_outputs(2786)));
    layer2_outputs(3348) <= layer1_outputs(731);
    layer2_outputs(3349) <= layer1_outputs(9893);
    layer2_outputs(3350) <= layer1_outputs(8084);
    layer2_outputs(3351) <= not((layer1_outputs(5430)) and (layer1_outputs(5370)));
    layer2_outputs(3352) <= (layer1_outputs(362)) and not (layer1_outputs(6312));
    layer2_outputs(3353) <= not(layer1_outputs(8603)) or (layer1_outputs(164));
    layer2_outputs(3354) <= not(layer1_outputs(8117));
    layer2_outputs(3355) <= not(layer1_outputs(7624));
    layer2_outputs(3356) <= layer1_outputs(9622);
    layer2_outputs(3357) <= layer1_outputs(1702);
    layer2_outputs(3358) <= not(layer1_outputs(7620)) or (layer1_outputs(8778));
    layer2_outputs(3359) <= layer1_outputs(7255);
    layer2_outputs(3360) <= not((layer1_outputs(4774)) and (layer1_outputs(1422)));
    layer2_outputs(3361) <= not((layer1_outputs(8251)) xor (layer1_outputs(3301)));
    layer2_outputs(3362) <= (layer1_outputs(7738)) and not (layer1_outputs(2080));
    layer2_outputs(3363) <= not(layer1_outputs(7798)) or (layer1_outputs(5645));
    layer2_outputs(3364) <= (layer1_outputs(8870)) and (layer1_outputs(9003));
    layer2_outputs(3365) <= layer1_outputs(8936);
    layer2_outputs(3366) <= layer1_outputs(3472);
    layer2_outputs(3367) <= layer1_outputs(5198);
    layer2_outputs(3368) <= layer1_outputs(4452);
    layer2_outputs(3369) <= not(layer1_outputs(9210));
    layer2_outputs(3370) <= layer1_outputs(4621);
    layer2_outputs(3371) <= layer1_outputs(469);
    layer2_outputs(3372) <= not((layer1_outputs(5860)) or (layer1_outputs(4089)));
    layer2_outputs(3373) <= not((layer1_outputs(6039)) or (layer1_outputs(5708)));
    layer2_outputs(3374) <= (layer1_outputs(7119)) xor (layer1_outputs(5890));
    layer2_outputs(3375) <= not(layer1_outputs(1131)) or (layer1_outputs(2035));
    layer2_outputs(3376) <= (layer1_outputs(9036)) xor (layer1_outputs(4794));
    layer2_outputs(3377) <= not(layer1_outputs(1710));
    layer2_outputs(3378) <= (layer1_outputs(7212)) xor (layer1_outputs(4524));
    layer2_outputs(3379) <= not(layer1_outputs(3839));
    layer2_outputs(3380) <= (layer1_outputs(2505)) and not (layer1_outputs(8531));
    layer2_outputs(3381) <= (layer1_outputs(3138)) and not (layer1_outputs(423));
    layer2_outputs(3382) <= not((layer1_outputs(346)) xor (layer1_outputs(8002)));
    layer2_outputs(3383) <= (layer1_outputs(5039)) and not (layer1_outputs(1879));
    layer2_outputs(3384) <= not(layer1_outputs(9927)) or (layer1_outputs(9022));
    layer2_outputs(3385) <= (layer1_outputs(4007)) and not (layer1_outputs(521));
    layer2_outputs(3386) <= layer1_outputs(9686);
    layer2_outputs(3387) <= layer1_outputs(815);
    layer2_outputs(3388) <= (layer1_outputs(2489)) xor (layer1_outputs(1034));
    layer2_outputs(3389) <= layer1_outputs(8402);
    layer2_outputs(3390) <= not((layer1_outputs(4513)) xor (layer1_outputs(4148)));
    layer2_outputs(3391) <= not(layer1_outputs(2194)) or (layer1_outputs(2283));
    layer2_outputs(3392) <= not(layer1_outputs(8679));
    layer2_outputs(3393) <= not(layer1_outputs(4035)) or (layer1_outputs(2069));
    layer2_outputs(3394) <= not(layer1_outputs(1779)) or (layer1_outputs(10014));
    layer2_outputs(3395) <= not(layer1_outputs(1921));
    layer2_outputs(3396) <= (layer1_outputs(1209)) or (layer1_outputs(7423));
    layer2_outputs(3397) <= (layer1_outputs(6922)) and not (layer1_outputs(2074));
    layer2_outputs(3398) <= not(layer1_outputs(3947));
    layer2_outputs(3399) <= (layer1_outputs(7428)) xor (layer1_outputs(6906));
    layer2_outputs(3400) <= (layer1_outputs(512)) xor (layer1_outputs(3171));
    layer2_outputs(3401) <= layer1_outputs(4283);
    layer2_outputs(3402) <= layer1_outputs(832);
    layer2_outputs(3403) <= layer1_outputs(303);
    layer2_outputs(3404) <= not(layer1_outputs(3880));
    layer2_outputs(3405) <= (layer1_outputs(8035)) and (layer1_outputs(5289));
    layer2_outputs(3406) <= layer1_outputs(7601);
    layer2_outputs(3407) <= not((layer1_outputs(1942)) xor (layer1_outputs(4414)));
    layer2_outputs(3408) <= layer1_outputs(7041);
    layer2_outputs(3409) <= layer1_outputs(1088);
    layer2_outputs(3410) <= not((layer1_outputs(5888)) and (layer1_outputs(3035)));
    layer2_outputs(3411) <= (layer1_outputs(4657)) and not (layer1_outputs(3733));
    layer2_outputs(3412) <= not((layer1_outputs(1372)) and (layer1_outputs(257)));
    layer2_outputs(3413) <= (layer1_outputs(3975)) or (layer1_outputs(1903));
    layer2_outputs(3414) <= not((layer1_outputs(3452)) xor (layer1_outputs(6581)));
    layer2_outputs(3415) <= not((layer1_outputs(285)) and (layer1_outputs(8528)));
    layer2_outputs(3416) <= layer1_outputs(7680);
    layer2_outputs(3417) <= layer1_outputs(9002);
    layer2_outputs(3418) <= (layer1_outputs(1571)) or (layer1_outputs(10037));
    layer2_outputs(3419) <= not(layer1_outputs(1474)) or (layer1_outputs(2505));
    layer2_outputs(3420) <= not(layer1_outputs(1233));
    layer2_outputs(3421) <= not(layer1_outputs(5215)) or (layer1_outputs(9057));
    layer2_outputs(3422) <= layer1_outputs(2567);
    layer2_outputs(3423) <= (layer1_outputs(5295)) or (layer1_outputs(3167));
    layer2_outputs(3424) <= not((layer1_outputs(5687)) and (layer1_outputs(2736)));
    layer2_outputs(3425) <= (layer1_outputs(9553)) and not (layer1_outputs(3764));
    layer2_outputs(3426) <= not((layer1_outputs(8127)) or (layer1_outputs(538)));
    layer2_outputs(3427) <= not(layer1_outputs(7898)) or (layer1_outputs(5035));
    layer2_outputs(3428) <= not((layer1_outputs(5204)) and (layer1_outputs(1160)));
    layer2_outputs(3429) <= not(layer1_outputs(1436));
    layer2_outputs(3430) <= not((layer1_outputs(5856)) or (layer1_outputs(9108)));
    layer2_outputs(3431) <= not(layer1_outputs(4946));
    layer2_outputs(3432) <= not((layer1_outputs(5536)) xor (layer1_outputs(937)));
    layer2_outputs(3433) <= (layer1_outputs(4233)) and (layer1_outputs(3611));
    layer2_outputs(3434) <= not(layer1_outputs(6302));
    layer2_outputs(3435) <= not(layer1_outputs(9261));
    layer2_outputs(3436) <= not(layer1_outputs(9138)) or (layer1_outputs(5906));
    layer2_outputs(3437) <= (layer1_outputs(5964)) and (layer1_outputs(308));
    layer2_outputs(3438) <= (layer1_outputs(513)) xor (layer1_outputs(7850));
    layer2_outputs(3439) <= not(layer1_outputs(8608));
    layer2_outputs(3440) <= not(layer1_outputs(9899));
    layer2_outputs(3441) <= '1';
    layer2_outputs(3442) <= layer1_outputs(9644);
    layer2_outputs(3443) <= layer1_outputs(6929);
    layer2_outputs(3444) <= not(layer1_outputs(580));
    layer2_outputs(3445) <= not((layer1_outputs(2768)) and (layer1_outputs(4190)));
    layer2_outputs(3446) <= not((layer1_outputs(8471)) or (layer1_outputs(7791)));
    layer2_outputs(3447) <= not(layer1_outputs(5273));
    layer2_outputs(3448) <= not((layer1_outputs(6001)) and (layer1_outputs(9371)));
    layer2_outputs(3449) <= (layer1_outputs(9051)) and (layer1_outputs(5742));
    layer2_outputs(3450) <= not(layer1_outputs(1506)) or (layer1_outputs(250));
    layer2_outputs(3451) <= layer1_outputs(5766);
    layer2_outputs(3452) <= not(layer1_outputs(1550));
    layer2_outputs(3453) <= (layer1_outputs(6945)) xor (layer1_outputs(4366));
    layer2_outputs(3454) <= not(layer1_outputs(5912));
    layer2_outputs(3455) <= (layer1_outputs(6486)) and (layer1_outputs(9433));
    layer2_outputs(3456) <= (layer1_outputs(1992)) or (layer1_outputs(7797));
    layer2_outputs(3457) <= layer1_outputs(8461);
    layer2_outputs(3458) <= not(layer1_outputs(9902));
    layer2_outputs(3459) <= (layer1_outputs(7626)) xor (layer1_outputs(4945));
    layer2_outputs(3460) <= not(layer1_outputs(9447));
    layer2_outputs(3461) <= not((layer1_outputs(9527)) xor (layer1_outputs(696)));
    layer2_outputs(3462) <= (layer1_outputs(151)) and not (layer1_outputs(6467));
    layer2_outputs(3463) <= not(layer1_outputs(7222));
    layer2_outputs(3464) <= not(layer1_outputs(3556));
    layer2_outputs(3465) <= not(layer1_outputs(5837));
    layer2_outputs(3466) <= not(layer1_outputs(7775));
    layer2_outputs(3467) <= layer1_outputs(5893);
    layer2_outputs(3468) <= (layer1_outputs(5089)) and (layer1_outputs(9313));
    layer2_outputs(3469) <= not(layer1_outputs(9711));
    layer2_outputs(3470) <= not((layer1_outputs(5985)) or (layer1_outputs(5838)));
    layer2_outputs(3471) <= not(layer1_outputs(2739));
    layer2_outputs(3472) <= (layer1_outputs(9321)) xor (layer1_outputs(318));
    layer2_outputs(3473) <= (layer1_outputs(2233)) and not (layer1_outputs(816));
    layer2_outputs(3474) <= (layer1_outputs(10189)) xor (layer1_outputs(9723));
    layer2_outputs(3475) <= layer1_outputs(4201);
    layer2_outputs(3476) <= not(layer1_outputs(8686));
    layer2_outputs(3477) <= layer1_outputs(9206);
    layer2_outputs(3478) <= not((layer1_outputs(7816)) and (layer1_outputs(5694)));
    layer2_outputs(3479) <= not(layer1_outputs(5383));
    layer2_outputs(3480) <= (layer1_outputs(7964)) and not (layer1_outputs(5758));
    layer2_outputs(3481) <= not((layer1_outputs(4241)) or (layer1_outputs(8301)));
    layer2_outputs(3482) <= not(layer1_outputs(7636)) or (layer1_outputs(2793));
    layer2_outputs(3483) <= (layer1_outputs(481)) xor (layer1_outputs(6322));
    layer2_outputs(3484) <= not(layer1_outputs(1015));
    layer2_outputs(3485) <= layer1_outputs(9274);
    layer2_outputs(3486) <= not(layer1_outputs(9061)) or (layer1_outputs(8077));
    layer2_outputs(3487) <= not((layer1_outputs(6410)) xor (layer1_outputs(10132)));
    layer2_outputs(3488) <= not((layer1_outputs(1222)) xor (layer1_outputs(6101)));
    layer2_outputs(3489) <= not(layer1_outputs(1060));
    layer2_outputs(3490) <= (layer1_outputs(2771)) and not (layer1_outputs(8131));
    layer2_outputs(3491) <= not(layer1_outputs(4790));
    layer2_outputs(3492) <= not(layer1_outputs(9727));
    layer2_outputs(3493) <= (layer1_outputs(1904)) or (layer1_outputs(1134));
    layer2_outputs(3494) <= not(layer1_outputs(9056));
    layer2_outputs(3495) <= layer1_outputs(5545);
    layer2_outputs(3496) <= not(layer1_outputs(3899));
    layer2_outputs(3497) <= layer1_outputs(4886);
    layer2_outputs(3498) <= layer1_outputs(494);
    layer2_outputs(3499) <= not(layer1_outputs(4898));
    layer2_outputs(3500) <= layer1_outputs(8109);
    layer2_outputs(3501) <= not(layer1_outputs(8054));
    layer2_outputs(3502) <= (layer1_outputs(5905)) and (layer1_outputs(4834));
    layer2_outputs(3503) <= not((layer1_outputs(3632)) or (layer1_outputs(5231)));
    layer2_outputs(3504) <= not((layer1_outputs(8712)) and (layer1_outputs(6218)));
    layer2_outputs(3505) <= not(layer1_outputs(6371));
    layer2_outputs(3506) <= layer1_outputs(6313);
    layer2_outputs(3507) <= not(layer1_outputs(2542));
    layer2_outputs(3508) <= not((layer1_outputs(1075)) or (layer1_outputs(4171)));
    layer2_outputs(3509) <= not(layer1_outputs(7053));
    layer2_outputs(3510) <= not(layer1_outputs(7036));
    layer2_outputs(3511) <= layer1_outputs(6175);
    layer2_outputs(3512) <= (layer1_outputs(9760)) or (layer1_outputs(3539));
    layer2_outputs(3513) <= layer1_outputs(2549);
    layer2_outputs(3514) <= not(layer1_outputs(4915));
    layer2_outputs(3515) <= not((layer1_outputs(7629)) or (layer1_outputs(4302)));
    layer2_outputs(3516) <= (layer1_outputs(8750)) or (layer1_outputs(6798));
    layer2_outputs(3517) <= not(layer1_outputs(2892));
    layer2_outputs(3518) <= layer1_outputs(9618);
    layer2_outputs(3519) <= layer1_outputs(9026);
    layer2_outputs(3520) <= (layer1_outputs(2881)) xor (layer1_outputs(6377));
    layer2_outputs(3521) <= layer1_outputs(4144);
    layer2_outputs(3522) <= not(layer1_outputs(7716)) or (layer1_outputs(3870));
    layer2_outputs(3523) <= not(layer1_outputs(4569));
    layer2_outputs(3524) <= not(layer1_outputs(4156));
    layer2_outputs(3525) <= not(layer1_outputs(3320));
    layer2_outputs(3526) <= not(layer1_outputs(3687));
    layer2_outputs(3527) <= layer1_outputs(952);
    layer2_outputs(3528) <= not(layer1_outputs(8070));
    layer2_outputs(3529) <= not((layer1_outputs(8809)) xor (layer1_outputs(6323)));
    layer2_outputs(3530) <= layer1_outputs(7360);
    layer2_outputs(3531) <= not((layer1_outputs(5216)) xor (layer1_outputs(4358)));
    layer2_outputs(3532) <= layer1_outputs(4752);
    layer2_outputs(3533) <= (layer1_outputs(2827)) and not (layer1_outputs(9843));
    layer2_outputs(3534) <= not(layer1_outputs(4075)) or (layer1_outputs(3201));
    layer2_outputs(3535) <= not(layer1_outputs(6635));
    layer2_outputs(3536) <= layer1_outputs(3270);
    layer2_outputs(3537) <= not((layer1_outputs(6073)) xor (layer1_outputs(7877)));
    layer2_outputs(3538) <= (layer1_outputs(466)) and (layer1_outputs(4557));
    layer2_outputs(3539) <= not((layer1_outputs(6272)) xor (layer1_outputs(7346)));
    layer2_outputs(3540) <= not(layer1_outputs(6624));
    layer2_outputs(3541) <= not(layer1_outputs(1112));
    layer2_outputs(3542) <= not(layer1_outputs(2785));
    layer2_outputs(3543) <= not((layer1_outputs(2857)) xor (layer1_outputs(2804)));
    layer2_outputs(3544) <= layer1_outputs(5997);
    layer2_outputs(3545) <= not((layer1_outputs(5550)) xor (layer1_outputs(6649)));
    layer2_outputs(3546) <= layer1_outputs(3424);
    layer2_outputs(3547) <= not((layer1_outputs(7818)) and (layer1_outputs(4163)));
    layer2_outputs(3548) <= not(layer1_outputs(6944));
    layer2_outputs(3549) <= layer1_outputs(2064);
    layer2_outputs(3550) <= not(layer1_outputs(2860));
    layer2_outputs(3551) <= layer1_outputs(3176);
    layer2_outputs(3552) <= not(layer1_outputs(8011));
    layer2_outputs(3553) <= (layer1_outputs(9123)) xor (layer1_outputs(7841));
    layer2_outputs(3554) <= not(layer1_outputs(1388));
    layer2_outputs(3555) <= layer1_outputs(1706);
    layer2_outputs(3556) <= (layer1_outputs(2037)) xor (layer1_outputs(3597));
    layer2_outputs(3557) <= not(layer1_outputs(1842));
    layer2_outputs(3558) <= not((layer1_outputs(3904)) xor (layer1_outputs(9586)));
    layer2_outputs(3559) <= not(layer1_outputs(5396));
    layer2_outputs(3560) <= (layer1_outputs(5504)) and (layer1_outputs(4028));
    layer2_outputs(3561) <= not(layer1_outputs(3247));
    layer2_outputs(3562) <= (layer1_outputs(7089)) and not (layer1_outputs(5091));
    layer2_outputs(3563) <= not(layer1_outputs(7655));
    layer2_outputs(3564) <= layer1_outputs(9850);
    layer2_outputs(3565) <= (layer1_outputs(3134)) and not (layer1_outputs(1851));
    layer2_outputs(3566) <= not(layer1_outputs(5165));
    layer2_outputs(3567) <= layer1_outputs(4731);
    layer2_outputs(3568) <= not((layer1_outputs(3682)) and (layer1_outputs(7157)));
    layer2_outputs(3569) <= (layer1_outputs(720)) and (layer1_outputs(1193));
    layer2_outputs(3570) <= layer1_outputs(2983);
    layer2_outputs(3571) <= layer1_outputs(2647);
    layer2_outputs(3572) <= not(layer1_outputs(3401));
    layer2_outputs(3573) <= (layer1_outputs(2882)) and not (layer1_outputs(8317));
    layer2_outputs(3574) <= not(layer1_outputs(8625));
    layer2_outputs(3575) <= (layer1_outputs(8359)) xor (layer1_outputs(7274));
    layer2_outputs(3576) <= not(layer1_outputs(8228));
    layer2_outputs(3577) <= not(layer1_outputs(1463)) or (layer1_outputs(8510));
    layer2_outputs(3578) <= layer1_outputs(2803);
    layer2_outputs(3579) <= layer1_outputs(5404);
    layer2_outputs(3580) <= (layer1_outputs(3146)) and (layer1_outputs(1947));
    layer2_outputs(3581) <= layer1_outputs(1400);
    layer2_outputs(3582) <= not(layer1_outputs(8067));
    layer2_outputs(3583) <= not((layer1_outputs(2086)) and (layer1_outputs(8664)));
    layer2_outputs(3584) <= (layer1_outputs(1067)) or (layer1_outputs(2176));
    layer2_outputs(3585) <= layer1_outputs(418);
    layer2_outputs(3586) <= (layer1_outputs(9849)) xor (layer1_outputs(6536));
    layer2_outputs(3587) <= layer1_outputs(1396);
    layer2_outputs(3588) <= not((layer1_outputs(5350)) or (layer1_outputs(3455)));
    layer2_outputs(3589) <= (layer1_outputs(9863)) and not (layer1_outputs(1468));
    layer2_outputs(3590) <= (layer1_outputs(1288)) and not (layer1_outputs(7851));
    layer2_outputs(3591) <= layer1_outputs(8791);
    layer2_outputs(3592) <= (layer1_outputs(6273)) and (layer1_outputs(2029));
    layer2_outputs(3593) <= not((layer1_outputs(7648)) and (layer1_outputs(5951)));
    layer2_outputs(3594) <= layer1_outputs(1038);
    layer2_outputs(3595) <= (layer1_outputs(9679)) and not (layer1_outputs(4939));
    layer2_outputs(3596) <= (layer1_outputs(1438)) and (layer1_outputs(4884));
    layer2_outputs(3597) <= not((layer1_outputs(8701)) and (layer1_outputs(9385)));
    layer2_outputs(3598) <= not(layer1_outputs(556)) or (layer1_outputs(8485));
    layer2_outputs(3599) <= not(layer1_outputs(2460));
    layer2_outputs(3600) <= not(layer1_outputs(2553));
    layer2_outputs(3601) <= layer1_outputs(6571);
    layer2_outputs(3602) <= not(layer1_outputs(160)) or (layer1_outputs(7075));
    layer2_outputs(3603) <= (layer1_outputs(271)) and (layer1_outputs(4396));
    layer2_outputs(3604) <= not((layer1_outputs(7065)) xor (layer1_outputs(3425)));
    layer2_outputs(3605) <= layer1_outputs(65);
    layer2_outputs(3606) <= (layer1_outputs(5827)) and not (layer1_outputs(1723));
    layer2_outputs(3607) <= layer1_outputs(6590);
    layer2_outputs(3608) <= layer1_outputs(5690);
    layer2_outputs(3609) <= (layer1_outputs(9477)) and (layer1_outputs(1825));
    layer2_outputs(3610) <= not((layer1_outputs(1840)) xor (layer1_outputs(4437)));
    layer2_outputs(3611) <= (layer1_outputs(123)) xor (layer1_outputs(1761));
    layer2_outputs(3612) <= not((layer1_outputs(8777)) xor (layer1_outputs(10124)));
    layer2_outputs(3613) <= layer1_outputs(6188);
    layer2_outputs(3614) <= layer1_outputs(4695);
    layer2_outputs(3615) <= (layer1_outputs(8389)) and not (layer1_outputs(10076));
    layer2_outputs(3616) <= layer1_outputs(855);
    layer2_outputs(3617) <= layer1_outputs(6316);
    layer2_outputs(3618) <= (layer1_outputs(7367)) xor (layer1_outputs(4574));
    layer2_outputs(3619) <= layer1_outputs(6925);
    layer2_outputs(3620) <= not((layer1_outputs(1175)) xor (layer1_outputs(1258)));
    layer2_outputs(3621) <= not(layer1_outputs(325)) or (layer1_outputs(6604));
    layer2_outputs(3622) <= not((layer1_outputs(7169)) or (layer1_outputs(1996)));
    layer2_outputs(3623) <= not(layer1_outputs(1822));
    layer2_outputs(3624) <= not(layer1_outputs(7270)) or (layer1_outputs(9517));
    layer2_outputs(3625) <= not(layer1_outputs(2349));
    layer2_outputs(3626) <= not(layer1_outputs(6666)) or (layer1_outputs(566));
    layer2_outputs(3627) <= layer1_outputs(2457);
    layer2_outputs(3628) <= layer1_outputs(7422);
    layer2_outputs(3629) <= layer1_outputs(9202);
    layer2_outputs(3630) <= layer1_outputs(2703);
    layer2_outputs(3631) <= not((layer1_outputs(2741)) xor (layer1_outputs(4567)));
    layer2_outputs(3632) <= layer1_outputs(402);
    layer2_outputs(3633) <= (layer1_outputs(10044)) xor (layer1_outputs(9884));
    layer2_outputs(3634) <= not(layer1_outputs(282));
    layer2_outputs(3635) <= (layer1_outputs(288)) or (layer1_outputs(2119));
    layer2_outputs(3636) <= layer1_outputs(9196);
    layer2_outputs(3637) <= layer1_outputs(6319);
    layer2_outputs(3638) <= layer1_outputs(8774);
    layer2_outputs(3639) <= not((layer1_outputs(6623)) xor (layer1_outputs(2765)));
    layer2_outputs(3640) <= layer1_outputs(7379);
    layer2_outputs(3641) <= layer1_outputs(986);
    layer2_outputs(3642) <= not(layer1_outputs(5740));
    layer2_outputs(3643) <= layer1_outputs(1235);
    layer2_outputs(3644) <= not(layer1_outputs(10062));
    layer2_outputs(3645) <= not(layer1_outputs(7729));
    layer2_outputs(3646) <= not((layer1_outputs(8439)) xor (layer1_outputs(351)));
    layer2_outputs(3647) <= not(layer1_outputs(7438));
    layer2_outputs(3648) <= not((layer1_outputs(654)) and (layer1_outputs(6193)));
    layer2_outputs(3649) <= not(layer1_outputs(5809));
    layer2_outputs(3650) <= not(layer1_outputs(2435));
    layer2_outputs(3651) <= layer1_outputs(6230);
    layer2_outputs(3652) <= not((layer1_outputs(7884)) or (layer1_outputs(9021)));
    layer2_outputs(3653) <= not(layer1_outputs(820));
    layer2_outputs(3654) <= not(layer1_outputs(2515));
    layer2_outputs(3655) <= layer1_outputs(6846);
    layer2_outputs(3656) <= layer1_outputs(2778);
    layer2_outputs(3657) <= layer1_outputs(9522);
    layer2_outputs(3658) <= not(layer1_outputs(10024)) or (layer1_outputs(6992));
    layer2_outputs(3659) <= not(layer1_outputs(2827)) or (layer1_outputs(9576));
    layer2_outputs(3660) <= not((layer1_outputs(3638)) xor (layer1_outputs(755)));
    layer2_outputs(3661) <= layer1_outputs(4583);
    layer2_outputs(3662) <= not((layer1_outputs(8007)) and (layer1_outputs(4538)));
    layer2_outputs(3663) <= (layer1_outputs(8852)) and not (layer1_outputs(5765));
    layer2_outputs(3664) <= not(layer1_outputs(627)) or (layer1_outputs(6175));
    layer2_outputs(3665) <= (layer1_outputs(314)) and (layer1_outputs(2426));
    layer2_outputs(3666) <= not(layer1_outputs(8710));
    layer2_outputs(3667) <= not(layer1_outputs(3959)) or (layer1_outputs(3587));
    layer2_outputs(3668) <= layer1_outputs(8905);
    layer2_outputs(3669) <= (layer1_outputs(3822)) and not (layer1_outputs(7565));
    layer2_outputs(3670) <= not(layer1_outputs(6555));
    layer2_outputs(3671) <= (layer1_outputs(9274)) and (layer1_outputs(2856));
    layer2_outputs(3672) <= (layer1_outputs(1894)) or (layer1_outputs(3447));
    layer2_outputs(3673) <= (layer1_outputs(6938)) and not (layer1_outputs(2196));
    layer2_outputs(3674) <= layer1_outputs(6667);
    layer2_outputs(3675) <= not((layer1_outputs(8568)) and (layer1_outputs(6094)));
    layer2_outputs(3676) <= not(layer1_outputs(8500));
    layer2_outputs(3677) <= not(layer1_outputs(2091)) or (layer1_outputs(9413));
    layer2_outputs(3678) <= not((layer1_outputs(5931)) xor (layer1_outputs(5512)));
    layer2_outputs(3679) <= not((layer1_outputs(10214)) or (layer1_outputs(6409)));
    layer2_outputs(3680) <= not(layer1_outputs(5756));
    layer2_outputs(3681) <= not(layer1_outputs(4420));
    layer2_outputs(3682) <= (layer1_outputs(4897)) xor (layer1_outputs(2177));
    layer2_outputs(3683) <= not((layer1_outputs(3841)) or (layer1_outputs(10020)));
    layer2_outputs(3684) <= not(layer1_outputs(397)) or (layer1_outputs(2955));
    layer2_outputs(3685) <= (layer1_outputs(5981)) and not (layer1_outputs(9645));
    layer2_outputs(3686) <= layer1_outputs(6840);
    layer2_outputs(3687) <= not((layer1_outputs(8672)) or (layer1_outputs(3344)));
    layer2_outputs(3688) <= layer1_outputs(7992);
    layer2_outputs(3689) <= not(layer1_outputs(3779)) or (layer1_outputs(6815));
    layer2_outputs(3690) <= layer1_outputs(8918);
    layer2_outputs(3691) <= not(layer1_outputs(4230));
    layer2_outputs(3692) <= not((layer1_outputs(7371)) or (layer1_outputs(3010)));
    layer2_outputs(3693) <= not((layer1_outputs(9001)) xor (layer1_outputs(1289)));
    layer2_outputs(3694) <= layer1_outputs(3091);
    layer2_outputs(3695) <= not(layer1_outputs(3903));
    layer2_outputs(3696) <= not((layer1_outputs(3678)) xor (layer1_outputs(2598)));
    layer2_outputs(3697) <= (layer1_outputs(5311)) and not (layer1_outputs(4144));
    layer2_outputs(3698) <= (layer1_outputs(3662)) and not (layer1_outputs(759));
    layer2_outputs(3699) <= not(layer1_outputs(6288));
    layer2_outputs(3700) <= not(layer1_outputs(5145)) or (layer1_outputs(12));
    layer2_outputs(3701) <= not(layer1_outputs(7699));
    layer2_outputs(3702) <= (layer1_outputs(6892)) or (layer1_outputs(5303));
    layer2_outputs(3703) <= not(layer1_outputs(558));
    layer2_outputs(3704) <= (layer1_outputs(2376)) and not (layer1_outputs(4598));
    layer2_outputs(3705) <= not((layer1_outputs(8307)) xor (layer1_outputs(1695)));
    layer2_outputs(3706) <= not(layer1_outputs(2097));
    layer2_outputs(3707) <= layer1_outputs(3665);
    layer2_outputs(3708) <= not(layer1_outputs(7514)) or (layer1_outputs(1521));
    layer2_outputs(3709) <= not(layer1_outputs(3490));
    layer2_outputs(3710) <= layer1_outputs(5203);
    layer2_outputs(3711) <= not((layer1_outputs(1483)) xor (layer1_outputs(2240)));
    layer2_outputs(3712) <= not(layer1_outputs(7276));
    layer2_outputs(3713) <= (layer1_outputs(9122)) or (layer1_outputs(5370));
    layer2_outputs(3714) <= not(layer1_outputs(7370));
    layer2_outputs(3715) <= not(layer1_outputs(5466));
    layer2_outputs(3716) <= not(layer1_outputs(873));
    layer2_outputs(3717) <= not((layer1_outputs(3924)) and (layer1_outputs(10099)));
    layer2_outputs(3718) <= not(layer1_outputs(5351));
    layer2_outputs(3719) <= not((layer1_outputs(5571)) xor (layer1_outputs(1736)));
    layer2_outputs(3720) <= (layer1_outputs(7210)) or (layer1_outputs(2622));
    layer2_outputs(3721) <= not((layer1_outputs(2451)) or (layer1_outputs(3791)));
    layer2_outputs(3722) <= layer1_outputs(7528);
    layer2_outputs(3723) <= layer1_outputs(3131);
    layer2_outputs(3724) <= not(layer1_outputs(646));
    layer2_outputs(3725) <= not(layer1_outputs(9078));
    layer2_outputs(3726) <= not((layer1_outputs(8794)) xor (layer1_outputs(2160)));
    layer2_outputs(3727) <= (layer1_outputs(3473)) or (layer1_outputs(9233));
    layer2_outputs(3728) <= not(layer1_outputs(3587));
    layer2_outputs(3729) <= not((layer1_outputs(3357)) or (layer1_outputs(2873)));
    layer2_outputs(3730) <= (layer1_outputs(7305)) and not (layer1_outputs(3030));
    layer2_outputs(3731) <= not(layer1_outputs(8528));
    layer2_outputs(3732) <= layer1_outputs(4887);
    layer2_outputs(3733) <= layer1_outputs(3372);
    layer2_outputs(3734) <= layer1_outputs(3683);
    layer2_outputs(3735) <= layer1_outputs(5168);
    layer2_outputs(3736) <= (layer1_outputs(4518)) and not (layer1_outputs(8838));
    layer2_outputs(3737) <= not((layer1_outputs(9334)) or (layer1_outputs(4770)));
    layer2_outputs(3738) <= not(layer1_outputs(7242));
    layer2_outputs(3739) <= (layer1_outputs(2912)) and not (layer1_outputs(8176));
    layer2_outputs(3740) <= not(layer1_outputs(8648)) or (layer1_outputs(5450));
    layer2_outputs(3741) <= (layer1_outputs(9272)) or (layer1_outputs(9573));
    layer2_outputs(3742) <= not(layer1_outputs(4140));
    layer2_outputs(3743) <= not(layer1_outputs(2314)) or (layer1_outputs(2396));
    layer2_outputs(3744) <= not(layer1_outputs(8147));
    layer2_outputs(3745) <= (layer1_outputs(4450)) xor (layer1_outputs(2287));
    layer2_outputs(3746) <= (layer1_outputs(3492)) and not (layer1_outputs(9888));
    layer2_outputs(3747) <= (layer1_outputs(234)) and not (layer1_outputs(4748));
    layer2_outputs(3748) <= not(layer1_outputs(3623));
    layer2_outputs(3749) <= not((layer1_outputs(452)) or (layer1_outputs(9488)));
    layer2_outputs(3750) <= layer1_outputs(7680);
    layer2_outputs(3751) <= layer1_outputs(5389);
    layer2_outputs(3752) <= not((layer1_outputs(1890)) xor (layer1_outputs(2779)));
    layer2_outputs(3753) <= not((layer1_outputs(3395)) or (layer1_outputs(9010)));
    layer2_outputs(3754) <= not(layer1_outputs(5969)) or (layer1_outputs(9875));
    layer2_outputs(3755) <= (layer1_outputs(1853)) and not (layer1_outputs(5638));
    layer2_outputs(3756) <= layer1_outputs(5319);
    layer2_outputs(3757) <= layer1_outputs(9103);
    layer2_outputs(3758) <= (layer1_outputs(4685)) xor (layer1_outputs(9084));
    layer2_outputs(3759) <= not((layer1_outputs(2471)) xor (layer1_outputs(8538)));
    layer2_outputs(3760) <= (layer1_outputs(2450)) and (layer1_outputs(4393));
    layer2_outputs(3761) <= not((layer1_outputs(1796)) or (layer1_outputs(10236)));
    layer2_outputs(3762) <= (layer1_outputs(2529)) and not (layer1_outputs(933));
    layer2_outputs(3763) <= not(layer1_outputs(6010)) or (layer1_outputs(3729));
    layer2_outputs(3764) <= layer1_outputs(5764);
    layer2_outputs(3765) <= not(layer1_outputs(7633));
    layer2_outputs(3766) <= not((layer1_outputs(5348)) and (layer1_outputs(6294)));
    layer2_outputs(3767) <= not(layer1_outputs(9737)) or (layer1_outputs(7385));
    layer2_outputs(3768) <= layer1_outputs(7670);
    layer2_outputs(3769) <= layer1_outputs(566);
    layer2_outputs(3770) <= (layer1_outputs(366)) and (layer1_outputs(4281));
    layer2_outputs(3771) <= not(layer1_outputs(8131));
    layer2_outputs(3772) <= (layer1_outputs(2178)) xor (layer1_outputs(3180));
    layer2_outputs(3773) <= not((layer1_outputs(4483)) or (layer1_outputs(653)));
    layer2_outputs(3774) <= layer1_outputs(623);
    layer2_outputs(3775) <= not(layer1_outputs(5334));
    layer2_outputs(3776) <= not(layer1_outputs(4334));
    layer2_outputs(3777) <= not((layer1_outputs(5477)) xor (layer1_outputs(623)));
    layer2_outputs(3778) <= not(layer1_outputs(5961));
    layer2_outputs(3779) <= (layer1_outputs(1640)) xor (layer1_outputs(6078));
    layer2_outputs(3780) <= (layer1_outputs(4473)) or (layer1_outputs(830));
    layer2_outputs(3781) <= layer1_outputs(377);
    layer2_outputs(3782) <= not((layer1_outputs(61)) and (layer1_outputs(7393)));
    layer2_outputs(3783) <= layer1_outputs(81);
    layer2_outputs(3784) <= (layer1_outputs(1532)) or (layer1_outputs(4841));
    layer2_outputs(3785) <= (layer1_outputs(10097)) or (layer1_outputs(4196));
    layer2_outputs(3786) <= not(layer1_outputs(713)) or (layer1_outputs(2158));
    layer2_outputs(3787) <= not((layer1_outputs(5218)) or (layer1_outputs(6530)));
    layer2_outputs(3788) <= (layer1_outputs(7667)) and not (layer1_outputs(5683));
    layer2_outputs(3789) <= not((layer1_outputs(7498)) xor (layer1_outputs(2102)));
    layer2_outputs(3790) <= layer1_outputs(3230);
    layer2_outputs(3791) <= not(layer1_outputs(8647));
    layer2_outputs(3792) <= not((layer1_outputs(9517)) xor (layer1_outputs(9124)));
    layer2_outputs(3793) <= layer1_outputs(7044);
    layer2_outputs(3794) <= (layer1_outputs(10222)) and not (layer1_outputs(5836));
    layer2_outputs(3795) <= layer1_outputs(5408);
    layer2_outputs(3796) <= not(layer1_outputs(1702));
    layer2_outputs(3797) <= not((layer1_outputs(1652)) xor (layer1_outputs(288)));
    layer2_outputs(3798) <= not(layer1_outputs(7435)) or (layer1_outputs(6277));
    layer2_outputs(3799) <= not(layer1_outputs(8123));
    layer2_outputs(3800) <= (layer1_outputs(4963)) and (layer1_outputs(942));
    layer2_outputs(3801) <= layer1_outputs(3199);
    layer2_outputs(3802) <= not(layer1_outputs(6384));
    layer2_outputs(3803) <= not((layer1_outputs(9840)) xor (layer1_outputs(7190)));
    layer2_outputs(3804) <= not((layer1_outputs(1527)) and (layer1_outputs(8153)));
    layer2_outputs(3805) <= not(layer1_outputs(7517));
    layer2_outputs(3806) <= not(layer1_outputs(2326)) or (layer1_outputs(8094));
    layer2_outputs(3807) <= layer1_outputs(2508);
    layer2_outputs(3808) <= (layer1_outputs(5178)) and (layer1_outputs(6557));
    layer2_outputs(3809) <= layer1_outputs(2195);
    layer2_outputs(3810) <= layer1_outputs(4064);
    layer2_outputs(3811) <= layer1_outputs(5268);
    layer2_outputs(3812) <= not(layer1_outputs(7559));
    layer2_outputs(3813) <= not(layer1_outputs(686));
    layer2_outputs(3814) <= (layer1_outputs(4909)) and (layer1_outputs(2750));
    layer2_outputs(3815) <= not(layer1_outputs(1169)) or (layer1_outputs(1389));
    layer2_outputs(3816) <= (layer1_outputs(4237)) or (layer1_outputs(4305));
    layer2_outputs(3817) <= not(layer1_outputs(15)) or (layer1_outputs(9328));
    layer2_outputs(3818) <= layer1_outputs(3750);
    layer2_outputs(3819) <= (layer1_outputs(2030)) and not (layer1_outputs(4265));
    layer2_outputs(3820) <= (layer1_outputs(8920)) and not (layer1_outputs(9052));
    layer2_outputs(3821) <= layer1_outputs(4827);
    layer2_outputs(3822) <= not(layer1_outputs(6825)) or (layer1_outputs(468));
    layer2_outputs(3823) <= (layer1_outputs(3796)) and not (layer1_outputs(6465));
    layer2_outputs(3824) <= (layer1_outputs(6997)) xor (layer1_outputs(1778));
    layer2_outputs(3825) <= not((layer1_outputs(1029)) xor (layer1_outputs(4677)));
    layer2_outputs(3826) <= layer1_outputs(7257);
    layer2_outputs(3827) <= (layer1_outputs(8003)) xor (layer1_outputs(1237));
    layer2_outputs(3828) <= (layer1_outputs(1401)) or (layer1_outputs(26));
    layer2_outputs(3829) <= not(layer1_outputs(626));
    layer2_outputs(3830) <= not((layer1_outputs(7970)) or (layer1_outputs(385)));
    layer2_outputs(3831) <= (layer1_outputs(2380)) and not (layer1_outputs(2257));
    layer2_outputs(3832) <= not((layer1_outputs(3717)) and (layer1_outputs(7468)));
    layer2_outputs(3833) <= (layer1_outputs(5190)) and not (layer1_outputs(6668));
    layer2_outputs(3834) <= not(layer1_outputs(8143));
    layer2_outputs(3835) <= layer1_outputs(4052);
    layer2_outputs(3836) <= layer1_outputs(2743);
    layer2_outputs(3837) <= not(layer1_outputs(2365)) or (layer1_outputs(4661));
    layer2_outputs(3838) <= layer1_outputs(9204);
    layer2_outputs(3839) <= (layer1_outputs(7183)) and not (layer1_outputs(8772));
    layer2_outputs(3840) <= (layer1_outputs(7572)) xor (layer1_outputs(10173));
    layer2_outputs(3841) <= not(layer1_outputs(6170)) or (layer1_outputs(1384));
    layer2_outputs(3842) <= layer1_outputs(8501);
    layer2_outputs(3843) <= (layer1_outputs(2386)) and not (layer1_outputs(4046));
    layer2_outputs(3844) <= not(layer1_outputs(5490)) or (layer1_outputs(582));
    layer2_outputs(3845) <= not(layer1_outputs(6064)) or (layer1_outputs(6381));
    layer2_outputs(3846) <= not(layer1_outputs(3697));
    layer2_outputs(3847) <= not((layer1_outputs(8848)) or (layer1_outputs(9778)));
    layer2_outputs(3848) <= (layer1_outputs(9898)) and (layer1_outputs(1352));
    layer2_outputs(3849) <= not(layer1_outputs(7356));
    layer2_outputs(3850) <= layer1_outputs(799);
    layer2_outputs(3851) <= not(layer1_outputs(9391)) or (layer1_outputs(8957));
    layer2_outputs(3852) <= not(layer1_outputs(4353));
    layer2_outputs(3853) <= not(layer1_outputs(8381));
    layer2_outputs(3854) <= (layer1_outputs(8253)) and (layer1_outputs(191));
    layer2_outputs(3855) <= not((layer1_outputs(366)) xor (layer1_outputs(7031)));
    layer2_outputs(3856) <= not(layer1_outputs(2283));
    layer2_outputs(3857) <= not(layer1_outputs(9100));
    layer2_outputs(3858) <= (layer1_outputs(2422)) xor (layer1_outputs(266));
    layer2_outputs(3859) <= layer1_outputs(6362);
    layer2_outputs(3860) <= not((layer1_outputs(6184)) and (layer1_outputs(131)));
    layer2_outputs(3861) <= layer1_outputs(8054);
    layer2_outputs(3862) <= not((layer1_outputs(9633)) and (layer1_outputs(8451)));
    layer2_outputs(3863) <= not((layer1_outputs(77)) xor (layer1_outputs(2042)));
    layer2_outputs(3864) <= not(layer1_outputs(7673)) or (layer1_outputs(4545));
    layer2_outputs(3865) <= not(layer1_outputs(700));
    layer2_outputs(3866) <= layer1_outputs(9024);
    layer2_outputs(3867) <= not((layer1_outputs(7994)) and (layer1_outputs(8556)));
    layer2_outputs(3868) <= (layer1_outputs(1335)) and (layer1_outputs(2465));
    layer2_outputs(3869) <= (layer1_outputs(4522)) and (layer1_outputs(1693));
    layer2_outputs(3870) <= layer1_outputs(5137);
    layer2_outputs(3871) <= not(layer1_outputs(6029));
    layer2_outputs(3872) <= layer1_outputs(6752);
    layer2_outputs(3873) <= not((layer1_outputs(8771)) xor (layer1_outputs(7358)));
    layer2_outputs(3874) <= not(layer1_outputs(10106));
    layer2_outputs(3875) <= layer1_outputs(6023);
    layer2_outputs(3876) <= (layer1_outputs(8462)) and not (layer1_outputs(6907));
    layer2_outputs(3877) <= (layer1_outputs(4993)) and (layer1_outputs(4161));
    layer2_outputs(3878) <= not(layer1_outputs(5264)) or (layer1_outputs(7858));
    layer2_outputs(3879) <= not(layer1_outputs(1948)) or (layer1_outputs(1059));
    layer2_outputs(3880) <= not((layer1_outputs(5524)) xor (layer1_outputs(6651)));
    layer2_outputs(3881) <= not(layer1_outputs(2605)) or (layer1_outputs(2775));
    layer2_outputs(3882) <= (layer1_outputs(5647)) and not (layer1_outputs(8863));
    layer2_outputs(3883) <= not((layer1_outputs(9162)) xor (layer1_outputs(9943)));
    layer2_outputs(3884) <= layer1_outputs(6667);
    layer2_outputs(3885) <= (layer1_outputs(9045)) and (layer1_outputs(7945));
    layer2_outputs(3886) <= (layer1_outputs(8381)) or (layer1_outputs(10034));
    layer2_outputs(3887) <= layer1_outputs(3814);
    layer2_outputs(3888) <= layer1_outputs(6286);
    layer2_outputs(3889) <= layer1_outputs(9334);
    layer2_outputs(3890) <= layer1_outputs(1280);
    layer2_outputs(3891) <= (layer1_outputs(7152)) xor (layer1_outputs(8453));
    layer2_outputs(3892) <= (layer1_outputs(1084)) and not (layer1_outputs(7054));
    layer2_outputs(3893) <= layer1_outputs(7777);
    layer2_outputs(3894) <= not(layer1_outputs(2747));
    layer2_outputs(3895) <= not(layer1_outputs(5225));
    layer2_outputs(3896) <= layer1_outputs(5993);
    layer2_outputs(3897) <= (layer1_outputs(4342)) and not (layer1_outputs(3344));
    layer2_outputs(3898) <= (layer1_outputs(3241)) and not (layer1_outputs(3274));
    layer2_outputs(3899) <= layer1_outputs(274);
    layer2_outputs(3900) <= (layer1_outputs(2091)) and not (layer1_outputs(4480));
    layer2_outputs(3901) <= not((layer1_outputs(1135)) xor (layer1_outputs(9311)));
    layer2_outputs(3902) <= not((layer1_outputs(652)) and (layer1_outputs(2253)));
    layer2_outputs(3903) <= layer1_outputs(1093);
    layer2_outputs(3904) <= layer1_outputs(9474);
    layer2_outputs(3905) <= not(layer1_outputs(5096));
    layer2_outputs(3906) <= layer1_outputs(1661);
    layer2_outputs(3907) <= layer1_outputs(4373);
    layer2_outputs(3908) <= layer1_outputs(6519);
    layer2_outputs(3909) <= layer1_outputs(9297);
    layer2_outputs(3910) <= not(layer1_outputs(8885));
    layer2_outputs(3911) <= not(layer1_outputs(5595));
    layer2_outputs(3912) <= (layer1_outputs(2239)) or (layer1_outputs(6419));
    layer2_outputs(3913) <= (layer1_outputs(7785)) or (layer1_outputs(1026));
    layer2_outputs(3914) <= (layer1_outputs(3225)) xor (layer1_outputs(10081));
    layer2_outputs(3915) <= layer1_outputs(4879);
    layer2_outputs(3916) <= not(layer1_outputs(6933));
    layer2_outputs(3917) <= layer1_outputs(8535);
    layer2_outputs(3918) <= layer1_outputs(880);
    layer2_outputs(3919) <= not(layer1_outputs(5298));
    layer2_outputs(3920) <= (layer1_outputs(6662)) and (layer1_outputs(9113));
    layer2_outputs(3921) <= (layer1_outputs(3180)) xor (layer1_outputs(1105));
    layer2_outputs(3922) <= (layer1_outputs(6902)) and not (layer1_outputs(1210));
    layer2_outputs(3923) <= not((layer1_outputs(5152)) and (layer1_outputs(7092)));
    layer2_outputs(3924) <= (layer1_outputs(1162)) xor (layer1_outputs(588));
    layer2_outputs(3925) <= not(layer1_outputs(1399));
    layer2_outputs(3926) <= (layer1_outputs(4104)) or (layer1_outputs(9059));
    layer2_outputs(3927) <= not(layer1_outputs(3965));
    layer2_outputs(3928) <= not((layer1_outputs(7998)) xor (layer1_outputs(434)));
    layer2_outputs(3929) <= layer1_outputs(1930);
    layer2_outputs(3930) <= layer1_outputs(1720);
    layer2_outputs(3931) <= not((layer1_outputs(8347)) or (layer1_outputs(2971)));
    layer2_outputs(3932) <= not(layer1_outputs(10009));
    layer2_outputs(3933) <= '0';
    layer2_outputs(3934) <= not(layer1_outputs(6910));
    layer2_outputs(3935) <= (layer1_outputs(3735)) xor (layer1_outputs(6658));
    layer2_outputs(3936) <= layer1_outputs(1037);
    layer2_outputs(3937) <= layer1_outputs(7657);
    layer2_outputs(3938) <= layer1_outputs(816);
    layer2_outputs(3939) <= not((layer1_outputs(894)) and (layer1_outputs(8611)));
    layer2_outputs(3940) <= layer1_outputs(5256);
    layer2_outputs(3941) <= (layer1_outputs(1603)) or (layer1_outputs(833));
    layer2_outputs(3942) <= layer1_outputs(9712);
    layer2_outputs(3943) <= not(layer1_outputs(2050));
    layer2_outputs(3944) <= (layer1_outputs(6641)) xor (layer1_outputs(348));
    layer2_outputs(3945) <= layer1_outputs(3287);
    layer2_outputs(3946) <= layer1_outputs(9347);
    layer2_outputs(3947) <= layer1_outputs(3365);
    layer2_outputs(3948) <= not(layer1_outputs(8074)) or (layer1_outputs(1906));
    layer2_outputs(3949) <= not((layer1_outputs(8430)) or (layer1_outputs(9998)));
    layer2_outputs(3950) <= layer1_outputs(2418);
    layer2_outputs(3951) <= (layer1_outputs(6513)) xor (layer1_outputs(3174));
    layer2_outputs(3952) <= not(layer1_outputs(10108)) or (layer1_outputs(3954));
    layer2_outputs(3953) <= (layer1_outputs(2271)) xor (layer1_outputs(5134));
    layer2_outputs(3954) <= layer1_outputs(7776);
    layer2_outputs(3955) <= not((layer1_outputs(2618)) xor (layer1_outputs(9324)));
    layer2_outputs(3956) <= layer1_outputs(6232);
    layer2_outputs(3957) <= not(layer1_outputs(5675)) or (layer1_outputs(4775));
    layer2_outputs(3958) <= layer1_outputs(6015);
    layer2_outputs(3959) <= layer1_outputs(8786);
    layer2_outputs(3960) <= not(layer1_outputs(5183));
    layer2_outputs(3961) <= layer1_outputs(4057);
    layer2_outputs(3962) <= not(layer1_outputs(8238));
    layer2_outputs(3963) <= layer1_outputs(1853);
    layer2_outputs(3964) <= not((layer1_outputs(5426)) and (layer1_outputs(2067)));
    layer2_outputs(3965) <= (layer1_outputs(3067)) xor (layer1_outputs(7954));
    layer2_outputs(3966) <= not(layer1_outputs(5108));
    layer2_outputs(3967) <= (layer1_outputs(9567)) or (layer1_outputs(764));
    layer2_outputs(3968) <= (layer1_outputs(3324)) or (layer1_outputs(2403));
    layer2_outputs(3969) <= not((layer1_outputs(8926)) or (layer1_outputs(3154)));
    layer2_outputs(3970) <= not(layer1_outputs(9065));
    layer2_outputs(3971) <= layer1_outputs(4017);
    layer2_outputs(3972) <= layer1_outputs(9792);
    layer2_outputs(3973) <= (layer1_outputs(9673)) and not (layer1_outputs(5902));
    layer2_outputs(3974) <= layer1_outputs(1809);
    layer2_outputs(3975) <= layer1_outputs(3818);
    layer2_outputs(3976) <= '0';
    layer2_outputs(3977) <= not((layer1_outputs(3718)) and (layer1_outputs(3932)));
    layer2_outputs(3978) <= (layer1_outputs(7917)) and (layer1_outputs(8507));
    layer2_outputs(3979) <= (layer1_outputs(6626)) and (layer1_outputs(7024));
    layer2_outputs(3980) <= not(layer1_outputs(1356));
    layer2_outputs(3981) <= not((layer1_outputs(5774)) xor (layer1_outputs(4280)));
    layer2_outputs(3982) <= (layer1_outputs(8363)) xor (layer1_outputs(8464));
    layer2_outputs(3983) <= layer1_outputs(4490);
    layer2_outputs(3984) <= not((layer1_outputs(7505)) or (layer1_outputs(8809)));
    layer2_outputs(3985) <= (layer1_outputs(5705)) and not (layer1_outputs(5137));
    layer2_outputs(3986) <= not((layer1_outputs(1657)) xor (layer1_outputs(1445)));
    layer2_outputs(3987) <= (layer1_outputs(8023)) and not (layer1_outputs(2039));
    layer2_outputs(3988) <= not(layer1_outputs(113)) or (layer1_outputs(5113));
    layer2_outputs(3989) <= not(layer1_outputs(1766));
    layer2_outputs(3990) <= not(layer1_outputs(9007));
    layer2_outputs(3991) <= (layer1_outputs(5917)) xor (layer1_outputs(5674));
    layer2_outputs(3992) <= not(layer1_outputs(592));
    layer2_outputs(3993) <= not((layer1_outputs(2446)) and (layer1_outputs(4728)));
    layer2_outputs(3994) <= not(layer1_outputs(1076));
    layer2_outputs(3995) <= layer1_outputs(7155);
    layer2_outputs(3996) <= layer1_outputs(444);
    layer2_outputs(3997) <= layer1_outputs(10060);
    layer2_outputs(3998) <= not(layer1_outputs(5197));
    layer2_outputs(3999) <= not((layer1_outputs(1813)) or (layer1_outputs(1579)));
    layer2_outputs(4000) <= (layer1_outputs(5107)) xor (layer1_outputs(4347));
    layer2_outputs(4001) <= (layer1_outputs(6891)) and not (layer1_outputs(5726));
    layer2_outputs(4002) <= not(layer1_outputs(7940)) or (layer1_outputs(5154));
    layer2_outputs(4003) <= (layer1_outputs(9457)) xor (layer1_outputs(801));
    layer2_outputs(4004) <= (layer1_outputs(446)) and (layer1_outputs(3217));
    layer2_outputs(4005) <= (layer1_outputs(8041)) or (layer1_outputs(2765));
    layer2_outputs(4006) <= not((layer1_outputs(9282)) xor (layer1_outputs(3804)));
    layer2_outputs(4007) <= layer1_outputs(8642);
    layer2_outputs(4008) <= (layer1_outputs(3944)) and not (layer1_outputs(8000));
    layer2_outputs(4009) <= (layer1_outputs(1863)) xor (layer1_outputs(6955));
    layer2_outputs(4010) <= not((layer1_outputs(4563)) xor (layer1_outputs(2710)));
    layer2_outputs(4011) <= not(layer1_outputs(8547));
    layer2_outputs(4012) <= not(layer1_outputs(5883));
    layer2_outputs(4013) <= (layer1_outputs(2806)) and (layer1_outputs(2227));
    layer2_outputs(4014) <= layer1_outputs(9849);
    layer2_outputs(4015) <= not(layer1_outputs(8235)) or (layer1_outputs(6813));
    layer2_outputs(4016) <= not((layer1_outputs(713)) and (layer1_outputs(235)));
    layer2_outputs(4017) <= not(layer1_outputs(4031));
    layer2_outputs(4018) <= not(layer1_outputs(3404)) or (layer1_outputs(5830));
    layer2_outputs(4019) <= layer1_outputs(7163);
    layer2_outputs(4020) <= (layer1_outputs(7479)) and (layer1_outputs(7137));
    layer2_outputs(4021) <= layer1_outputs(6300);
    layer2_outputs(4022) <= not((layer1_outputs(8075)) xor (layer1_outputs(5824)));
    layer2_outputs(4023) <= not((layer1_outputs(10202)) and (layer1_outputs(9302)));
    layer2_outputs(4024) <= layer1_outputs(8289);
    layer2_outputs(4025) <= (layer1_outputs(3245)) xor (layer1_outputs(3760));
    layer2_outputs(4026) <= layer1_outputs(9343);
    layer2_outputs(4027) <= (layer1_outputs(1963)) and (layer1_outputs(9450));
    layer2_outputs(4028) <= not(layer1_outputs(1395));
    layer2_outputs(4029) <= (layer1_outputs(7590)) and not (layer1_outputs(10064));
    layer2_outputs(4030) <= layer1_outputs(1089);
    layer2_outputs(4031) <= (layer1_outputs(975)) and not (layer1_outputs(10220));
    layer2_outputs(4032) <= (layer1_outputs(6479)) and not (layer1_outputs(1600));
    layer2_outputs(4033) <= not(layer1_outputs(305));
    layer2_outputs(4034) <= (layer1_outputs(8969)) and not (layer1_outputs(9997));
    layer2_outputs(4035) <= layer1_outputs(214);
    layer2_outputs(4036) <= not((layer1_outputs(2733)) and (layer1_outputs(6140)));
    layer2_outputs(4037) <= not(layer1_outputs(3626)) or (layer1_outputs(9822));
    layer2_outputs(4038) <= not(layer1_outputs(6147)) or (layer1_outputs(9935));
    layer2_outputs(4039) <= not(layer1_outputs(6877));
    layer2_outputs(4040) <= not(layer1_outputs(6912)) or (layer1_outputs(6960));
    layer2_outputs(4041) <= (layer1_outputs(4701)) xor (layer1_outputs(8670));
    layer2_outputs(4042) <= layer1_outputs(4832);
    layer2_outputs(4043) <= not(layer1_outputs(3039));
    layer2_outputs(4044) <= not((layer1_outputs(9573)) or (layer1_outputs(7480)));
    layer2_outputs(4045) <= (layer1_outputs(9460)) xor (layer1_outputs(8696));
    layer2_outputs(4046) <= not((layer1_outputs(473)) xor (layer1_outputs(2181)));
    layer2_outputs(4047) <= layer1_outputs(9241);
    layer2_outputs(4048) <= not((layer1_outputs(10182)) xor (layer1_outputs(3560)));
    layer2_outputs(4049) <= not(layer1_outputs(3174));
    layer2_outputs(4050) <= not(layer1_outputs(373)) or (layer1_outputs(8407));
    layer2_outputs(4051) <= layer1_outputs(7763);
    layer2_outputs(4052) <= (layer1_outputs(1814)) or (layer1_outputs(1175));
    layer2_outputs(4053) <= (layer1_outputs(5679)) and not (layer1_outputs(538));
    layer2_outputs(4054) <= layer1_outputs(1950);
    layer2_outputs(4055) <= not(layer1_outputs(205));
    layer2_outputs(4056) <= not(layer1_outputs(5520));
    layer2_outputs(4057) <= layer1_outputs(7442);
    layer2_outputs(4058) <= not((layer1_outputs(9915)) and (layer1_outputs(4418)));
    layer2_outputs(4059) <= not(layer1_outputs(2697));
    layer2_outputs(4060) <= (layer1_outputs(5729)) and not (layer1_outputs(910));
    layer2_outputs(4061) <= layer1_outputs(210);
    layer2_outputs(4062) <= not(layer1_outputs(9598));
    layer2_outputs(4063) <= (layer1_outputs(1504)) xor (layer1_outputs(5146));
    layer2_outputs(4064) <= not(layer1_outputs(3275));
    layer2_outputs(4065) <= layer1_outputs(4361);
    layer2_outputs(4066) <= not((layer1_outputs(6014)) or (layer1_outputs(4717)));
    layer2_outputs(4067) <= not(layer1_outputs(8772));
    layer2_outputs(4068) <= (layer1_outputs(8910)) or (layer1_outputs(4639));
    layer2_outputs(4069) <= layer1_outputs(6743);
    layer2_outputs(4070) <= layer1_outputs(8355);
    layer2_outputs(4071) <= not(layer1_outputs(8638)) or (layer1_outputs(3545));
    layer2_outputs(4072) <= not(layer1_outputs(5076));
    layer2_outputs(4073) <= not((layer1_outputs(4577)) xor (layer1_outputs(2509)));
    layer2_outputs(4074) <= not(layer1_outputs(10112));
    layer2_outputs(4075) <= not((layer1_outputs(5872)) and (layer1_outputs(2235)));
    layer2_outputs(4076) <= not(layer1_outputs(6035));
    layer2_outputs(4077) <= not(layer1_outputs(2686));
    layer2_outputs(4078) <= (layer1_outputs(7805)) and (layer1_outputs(6363));
    layer2_outputs(4079) <= not(layer1_outputs(4103));
    layer2_outputs(4080) <= layer1_outputs(521);
    layer2_outputs(4081) <= '0';
    layer2_outputs(4082) <= layer1_outputs(9592);
    layer2_outputs(4083) <= not((layer1_outputs(8671)) and (layer1_outputs(4060)));
    layer2_outputs(4084) <= (layer1_outputs(1804)) or (layer1_outputs(4031));
    layer2_outputs(4085) <= not(layer1_outputs(6698));
    layer2_outputs(4086) <= not(layer1_outputs(606)) or (layer1_outputs(8261));
    layer2_outputs(4087) <= not((layer1_outputs(5541)) or (layer1_outputs(1006)));
    layer2_outputs(4088) <= (layer1_outputs(8220)) xor (layer1_outputs(6098));
    layer2_outputs(4089) <= not(layer1_outputs(6621)) or (layer1_outputs(3397));
    layer2_outputs(4090) <= (layer1_outputs(6499)) and not (layer1_outputs(8191));
    layer2_outputs(4091) <= layer1_outputs(2516);
    layer2_outputs(4092) <= not((layer1_outputs(7629)) xor (layer1_outputs(5330)));
    layer2_outputs(4093) <= layer1_outputs(6503);
    layer2_outputs(4094) <= not((layer1_outputs(3928)) or (layer1_outputs(5694)));
    layer2_outputs(4095) <= not(layer1_outputs(5543));
    layer2_outputs(4096) <= not(layer1_outputs(6449));
    layer2_outputs(4097) <= not(layer1_outputs(2731));
    layer2_outputs(4098) <= not(layer1_outputs(4203));
    layer2_outputs(4099) <= not(layer1_outputs(2188));
    layer2_outputs(4100) <= not(layer1_outputs(4462));
    layer2_outputs(4101) <= (layer1_outputs(2698)) and not (layer1_outputs(6519));
    layer2_outputs(4102) <= not(layer1_outputs(2520));
    layer2_outputs(4103) <= (layer1_outputs(3514)) or (layer1_outputs(10021));
    layer2_outputs(4104) <= not(layer1_outputs(7918));
    layer2_outputs(4105) <= (layer1_outputs(2705)) xor (layer1_outputs(6686));
    layer2_outputs(4106) <= not((layer1_outputs(5644)) or (layer1_outputs(3127)));
    layer2_outputs(4107) <= not(layer1_outputs(983)) or (layer1_outputs(8398));
    layer2_outputs(4108) <= (layer1_outputs(3330)) or (layer1_outputs(5034));
    layer2_outputs(4109) <= not(layer1_outputs(5772));
    layer2_outputs(4110) <= layer1_outputs(6020);
    layer2_outputs(4111) <= (layer1_outputs(7984)) and not (layer1_outputs(2288));
    layer2_outputs(4112) <= not(layer1_outputs(8516)) or (layer1_outputs(7392));
    layer2_outputs(4113) <= (layer1_outputs(4051)) and not (layer1_outputs(8453));
    layer2_outputs(4114) <= not(layer1_outputs(4636));
    layer2_outputs(4115) <= not((layer1_outputs(6151)) or (layer1_outputs(861)));
    layer2_outputs(4116) <= not(layer1_outputs(2078));
    layer2_outputs(4117) <= not((layer1_outputs(227)) or (layer1_outputs(4880)));
    layer2_outputs(4118) <= not(layer1_outputs(9705)) or (layer1_outputs(4));
    layer2_outputs(4119) <= layer1_outputs(842);
    layer2_outputs(4120) <= layer1_outputs(5783);
    layer2_outputs(4121) <= not(layer1_outputs(4760));
    layer2_outputs(4122) <= layer1_outputs(4377);
    layer2_outputs(4123) <= layer1_outputs(2830);
    layer2_outputs(4124) <= not(layer1_outputs(5387)) or (layer1_outputs(10141));
    layer2_outputs(4125) <= '0';
    layer2_outputs(4126) <= layer1_outputs(9384);
    layer2_outputs(4127) <= not(layer1_outputs(7308)) or (layer1_outputs(4374));
    layer2_outputs(4128) <= not(layer1_outputs(7814)) or (layer1_outputs(9441));
    layer2_outputs(4129) <= not(layer1_outputs(8277));
    layer2_outputs(4130) <= not((layer1_outputs(9025)) xor (layer1_outputs(8241)));
    layer2_outputs(4131) <= not(layer1_outputs(3738));
    layer2_outputs(4132) <= (layer1_outputs(9946)) and not (layer1_outputs(8742));
    layer2_outputs(4133) <= (layer1_outputs(1366)) and not (layer1_outputs(5274));
    layer2_outputs(4134) <= not(layer1_outputs(8928));
    layer2_outputs(4135) <= not((layer1_outputs(2852)) or (layer1_outputs(10190)));
    layer2_outputs(4136) <= not(layer1_outputs(2934)) or (layer1_outputs(4141));
    layer2_outputs(4137) <= (layer1_outputs(10158)) and not (layer1_outputs(6715));
    layer2_outputs(4138) <= layer1_outputs(5095);
    layer2_outputs(4139) <= not(layer1_outputs(8034)) or (layer1_outputs(7329));
    layer2_outputs(4140) <= not(layer1_outputs(1281));
    layer2_outputs(4141) <= not(layer1_outputs(4488));
    layer2_outputs(4142) <= not(layer1_outputs(3440)) or (layer1_outputs(8671));
    layer2_outputs(4143) <= not(layer1_outputs(3346));
    layer2_outputs(4144) <= (layer1_outputs(5158)) xor (layer1_outputs(3612));
    layer2_outputs(4145) <= (layer1_outputs(7673)) or (layer1_outputs(7766));
    layer2_outputs(4146) <= layer1_outputs(7148);
    layer2_outputs(4147) <= not(layer1_outputs(1124));
    layer2_outputs(4148) <= not(layer1_outputs(9701)) or (layer1_outputs(4867));
    layer2_outputs(4149) <= not(layer1_outputs(1440));
    layer2_outputs(4150) <= layer1_outputs(6535);
    layer2_outputs(4151) <= not(layer1_outputs(6252)) or (layer1_outputs(5298));
    layer2_outputs(4152) <= not(layer1_outputs(8272));
    layer2_outputs(4153) <= (layer1_outputs(4576)) xor (layer1_outputs(2183));
    layer2_outputs(4154) <= (layer1_outputs(9722)) xor (layer1_outputs(7081));
    layer2_outputs(4155) <= (layer1_outputs(3041)) and not (layer1_outputs(7050));
    layer2_outputs(4156) <= not((layer1_outputs(5790)) or (layer1_outputs(9908)));
    layer2_outputs(4157) <= (layer1_outputs(1104)) and not (layer1_outputs(2877));
    layer2_outputs(4158) <= layer1_outputs(6919);
    layer2_outputs(4159) <= not(layer1_outputs(3554)) or (layer1_outputs(6199));
    layer2_outputs(4160) <= layer1_outputs(8958);
    layer2_outputs(4161) <= (layer1_outputs(5288)) xor (layer1_outputs(2704));
    layer2_outputs(4162) <= not(layer1_outputs(2764));
    layer2_outputs(4163) <= not(layer1_outputs(2216)) or (layer1_outputs(8996));
    layer2_outputs(4164) <= not(layer1_outputs(4357));
    layer2_outputs(4165) <= not((layer1_outputs(8424)) and (layer1_outputs(6966)));
    layer2_outputs(4166) <= layer1_outputs(8323);
    layer2_outputs(4167) <= layer1_outputs(5813);
    layer2_outputs(4168) <= (layer1_outputs(3229)) xor (layer1_outputs(7790));
    layer2_outputs(4169) <= not((layer1_outputs(9820)) xor (layer1_outputs(2818)));
    layer2_outputs(4170) <= not(layer1_outputs(7145));
    layer2_outputs(4171) <= not(layer1_outputs(8329));
    layer2_outputs(4172) <= (layer1_outputs(1622)) and (layer1_outputs(7448));
    layer2_outputs(4173) <= not(layer1_outputs(9226)) or (layer1_outputs(6205));
    layer2_outputs(4174) <= (layer1_outputs(5724)) and not (layer1_outputs(6859));
    layer2_outputs(4175) <= not((layer1_outputs(3704)) xor (layer1_outputs(3412)));
    layer2_outputs(4176) <= not(layer1_outputs(8297)) or (layer1_outputs(311));
    layer2_outputs(4177) <= layer1_outputs(8256);
    layer2_outputs(4178) <= not(layer1_outputs(4225)) or (layer1_outputs(5501));
    layer2_outputs(4179) <= not((layer1_outputs(5795)) or (layer1_outputs(3928)));
    layer2_outputs(4180) <= not(layer1_outputs(6031));
    layer2_outputs(4181) <= layer1_outputs(8736);
    layer2_outputs(4182) <= not(layer1_outputs(9222));
    layer2_outputs(4183) <= not(layer1_outputs(10208));
    layer2_outputs(4184) <= not(layer1_outputs(6395));
    layer2_outputs(4185) <= (layer1_outputs(5294)) and not (layer1_outputs(4249));
    layer2_outputs(4186) <= not((layer1_outputs(2874)) or (layer1_outputs(3943)));
    layer2_outputs(4187) <= not(layer1_outputs(2494));
    layer2_outputs(4188) <= not(layer1_outputs(1503));
    layer2_outputs(4189) <= (layer1_outputs(5377)) xor (layer1_outputs(4217));
    layer2_outputs(4190) <= (layer1_outputs(6183)) and not (layer1_outputs(7304));
    layer2_outputs(4191) <= layer1_outputs(4381);
    layer2_outputs(4192) <= (layer1_outputs(2315)) xor (layer1_outputs(8829));
    layer2_outputs(4193) <= layer1_outputs(1441);
    layer2_outputs(4194) <= not((layer1_outputs(1927)) or (layer1_outputs(7076)));
    layer2_outputs(4195) <= (layer1_outputs(5429)) and (layer1_outputs(7264));
    layer2_outputs(4196) <= (layer1_outputs(2152)) xor (layer1_outputs(9040));
    layer2_outputs(4197) <= not((layer1_outputs(5121)) or (layer1_outputs(7292)));
    layer2_outputs(4198) <= (layer1_outputs(3212)) and (layer1_outputs(2024));
    layer2_outputs(4199) <= not(layer1_outputs(6755)) or (layer1_outputs(3526));
    layer2_outputs(4200) <= layer1_outputs(2036);
    layer2_outputs(4201) <= (layer1_outputs(7837)) xor (layer1_outputs(6765));
    layer2_outputs(4202) <= (layer1_outputs(10149)) and not (layer1_outputs(3118));
    layer2_outputs(4203) <= not(layer1_outputs(476));
    layer2_outputs(4204) <= not(layer1_outputs(2782));
    layer2_outputs(4205) <= not(layer1_outputs(5462)) or (layer1_outputs(2169));
    layer2_outputs(4206) <= (layer1_outputs(8185)) or (layer1_outputs(5839));
    layer2_outputs(4207) <= (layer1_outputs(8401)) and not (layer1_outputs(1574));
    layer2_outputs(4208) <= not((layer1_outputs(4019)) xor (layer1_outputs(4247)));
    layer2_outputs(4209) <= not(layer1_outputs(9150)) or (layer1_outputs(8562));
    layer2_outputs(4210) <= (layer1_outputs(8636)) xor (layer1_outputs(6154));
    layer2_outputs(4211) <= (layer1_outputs(3561)) and (layer1_outputs(3417));
    layer2_outputs(4212) <= layer1_outputs(5573);
    layer2_outputs(4213) <= layer1_outputs(8647);
    layer2_outputs(4214) <= layer1_outputs(6846);
    layer2_outputs(4215) <= layer1_outputs(5336);
    layer2_outputs(4216) <= (layer1_outputs(7604)) and not (layer1_outputs(1478));
    layer2_outputs(4217) <= layer1_outputs(10089);
    layer2_outputs(4218) <= not(layer1_outputs(4029));
    layer2_outputs(4219) <= layer1_outputs(6990);
    layer2_outputs(4220) <= (layer1_outputs(1781)) and not (layer1_outputs(1050));
    layer2_outputs(4221) <= layer1_outputs(7757);
    layer2_outputs(4222) <= '0';
    layer2_outputs(4223) <= not((layer1_outputs(1867)) and (layer1_outputs(5870)));
    layer2_outputs(4224) <= not(layer1_outputs(2565)) or (layer1_outputs(342));
    layer2_outputs(4225) <= layer1_outputs(496);
    layer2_outputs(4226) <= (layer1_outputs(7260)) or (layer1_outputs(3242));
    layer2_outputs(4227) <= not(layer1_outputs(2806)) or (layer1_outputs(58));
    layer2_outputs(4228) <= not(layer1_outputs(1808));
    layer2_outputs(4229) <= not(layer1_outputs(3938)) or (layer1_outputs(5010));
    layer2_outputs(4230) <= layer1_outputs(3252);
    layer2_outputs(4231) <= not((layer1_outputs(5181)) or (layer1_outputs(1951)));
    layer2_outputs(4232) <= not(layer1_outputs(7040));
    layer2_outputs(4233) <= (layer1_outputs(3021)) xor (layer1_outputs(9115));
    layer2_outputs(4234) <= not((layer1_outputs(9542)) xor (layer1_outputs(11)));
    layer2_outputs(4235) <= not(layer1_outputs(1506));
    layer2_outputs(4236) <= layer1_outputs(6339);
    layer2_outputs(4237) <= not(layer1_outputs(1164));
    layer2_outputs(4238) <= not((layer1_outputs(1042)) and (layer1_outputs(6775)));
    layer2_outputs(4239) <= layer1_outputs(9293);
    layer2_outputs(4240) <= not(layer1_outputs(4107));
    layer2_outputs(4241) <= not(layer1_outputs(8753));
    layer2_outputs(4242) <= not(layer1_outputs(3991));
    layer2_outputs(4243) <= layer1_outputs(8743);
    layer2_outputs(4244) <= (layer1_outputs(4453)) or (layer1_outputs(9497));
    layer2_outputs(4245) <= layer1_outputs(5792);
    layer2_outputs(4246) <= (layer1_outputs(9218)) xor (layer1_outputs(9527));
    layer2_outputs(4247) <= layer1_outputs(3639);
    layer2_outputs(4248) <= '1';
    layer2_outputs(4249) <= (layer1_outputs(6899)) and not (layer1_outputs(6931));
    layer2_outputs(4250) <= not(layer1_outputs(2713)) or (layer1_outputs(378));
    layer2_outputs(4251) <= not(layer1_outputs(9292)) or (layer1_outputs(5385));
    layer2_outputs(4252) <= (layer1_outputs(6332)) or (layer1_outputs(2142));
    layer2_outputs(4253) <= layer1_outputs(5367);
    layer2_outputs(4254) <= not(layer1_outputs(3973));
    layer2_outputs(4255) <= not(layer1_outputs(2600));
    layer2_outputs(4256) <= not((layer1_outputs(1377)) xor (layer1_outputs(4028)));
    layer2_outputs(4257) <= not(layer1_outputs(8722));
    layer2_outputs(4258) <= layer1_outputs(9550);
    layer2_outputs(4259) <= (layer1_outputs(10153)) and not (layer1_outputs(807));
    layer2_outputs(4260) <= (layer1_outputs(7310)) and (layer1_outputs(7269));
    layer2_outputs(4261) <= not(layer1_outputs(2381));
    layer2_outputs(4262) <= '0';
    layer2_outputs(4263) <= not(layer1_outputs(6732));
    layer2_outputs(4264) <= (layer1_outputs(4190)) xor (layer1_outputs(4402));
    layer2_outputs(4265) <= layer1_outputs(6946);
    layer2_outputs(4266) <= layer1_outputs(3551);
    layer2_outputs(4267) <= not(layer1_outputs(7682));
    layer2_outputs(4268) <= layer1_outputs(2957);
    layer2_outputs(4269) <= (layer1_outputs(7573)) and not (layer1_outputs(883));
    layer2_outputs(4270) <= not(layer1_outputs(7575));
    layer2_outputs(4271) <= not(layer1_outputs(6763));
    layer2_outputs(4272) <= layer1_outputs(8006);
    layer2_outputs(4273) <= not((layer1_outputs(2490)) xor (layer1_outputs(9199)));
    layer2_outputs(4274) <= (layer1_outputs(4276)) xor (layer1_outputs(3702));
    layer2_outputs(4275) <= (layer1_outputs(9317)) xor (layer1_outputs(7322));
    layer2_outputs(4276) <= not(layer1_outputs(3955));
    layer2_outputs(4277) <= not(layer1_outputs(5369));
    layer2_outputs(4278) <= not(layer1_outputs(5411));
    layer2_outputs(4279) <= not(layer1_outputs(5858)) or (layer1_outputs(9119));
    layer2_outputs(4280) <= not(layer1_outputs(10139));
    layer2_outputs(4281) <= (layer1_outputs(2766)) or (layer1_outputs(9271));
    layer2_outputs(4282) <= layer1_outputs(10227);
    layer2_outputs(4283) <= not((layer1_outputs(5702)) and (layer1_outputs(5432)));
    layer2_outputs(4284) <= (layer1_outputs(9995)) and not (layer1_outputs(6612));
    layer2_outputs(4285) <= (layer1_outputs(6053)) and not (layer1_outputs(7530));
    layer2_outputs(4286) <= (layer1_outputs(8612)) and (layer1_outputs(28));
    layer2_outputs(4287) <= (layer1_outputs(3218)) and not (layer1_outputs(5191));
    layer2_outputs(4288) <= (layer1_outputs(2959)) xor (layer1_outputs(8688));
    layer2_outputs(4289) <= layer1_outputs(638);
    layer2_outputs(4290) <= not(layer1_outputs(795));
    layer2_outputs(4291) <= not((layer1_outputs(7992)) or (layer1_outputs(174)));
    layer2_outputs(4292) <= not(layer1_outputs(7527));
    layer2_outputs(4293) <= not(layer1_outputs(10136));
    layer2_outputs(4294) <= not(layer1_outputs(7046)) or (layer1_outputs(9335));
    layer2_outputs(4295) <= not(layer1_outputs(8403));
    layer2_outputs(4296) <= not(layer1_outputs(5970));
    layer2_outputs(4297) <= (layer1_outputs(3388)) or (layer1_outputs(196));
    layer2_outputs(4298) <= not(layer1_outputs(3426)) or (layer1_outputs(472));
    layer2_outputs(4299) <= not(layer1_outputs(3478));
    layer2_outputs(4300) <= layer1_outputs(3393);
    layer2_outputs(4301) <= not(layer1_outputs(29)) or (layer1_outputs(3726));
    layer2_outputs(4302) <= (layer1_outputs(9837)) and (layer1_outputs(945));
    layer2_outputs(4303) <= not(layer1_outputs(6337));
    layer2_outputs(4304) <= not(layer1_outputs(7997)) or (layer1_outputs(1829));
    layer2_outputs(4305) <= not(layer1_outputs(5992)) or (layer1_outputs(7137));
    layer2_outputs(4306) <= not(layer1_outputs(1199));
    layer2_outputs(4307) <= not((layer1_outputs(5956)) or (layer1_outputs(908)));
    layer2_outputs(4308) <= not((layer1_outputs(3436)) and (layer1_outputs(8793)));
    layer2_outputs(4309) <= not(layer1_outputs(8050)) or (layer1_outputs(7849));
    layer2_outputs(4310) <= (layer1_outputs(1548)) and not (layer1_outputs(8146));
    layer2_outputs(4311) <= not(layer1_outputs(1173));
    layer2_outputs(4312) <= not(layer1_outputs(4147));
    layer2_outputs(4313) <= not(layer1_outputs(2643));
    layer2_outputs(4314) <= (layer1_outputs(2663)) and not (layer1_outputs(4625));
    layer2_outputs(4315) <= layer1_outputs(7043);
    layer2_outputs(4316) <= (layer1_outputs(2022)) and not (layer1_outputs(9044));
    layer2_outputs(4317) <= (layer1_outputs(10150)) xor (layer1_outputs(4375));
    layer2_outputs(4318) <= not((layer1_outputs(8856)) xor (layer1_outputs(9780)));
    layer2_outputs(4319) <= (layer1_outputs(8113)) and not (layer1_outputs(3189));
    layer2_outputs(4320) <= not(layer1_outputs(4549)) or (layer1_outputs(3614));
    layer2_outputs(4321) <= not(layer1_outputs(2610));
    layer2_outputs(4322) <= not(layer1_outputs(5465));
    layer2_outputs(4323) <= layer1_outputs(518);
    layer2_outputs(4324) <= not(layer1_outputs(863));
    layer2_outputs(4325) <= layer1_outputs(3541);
    layer2_outputs(4326) <= layer1_outputs(8442);
    layer2_outputs(4327) <= (layer1_outputs(14)) and not (layer1_outputs(7418));
    layer2_outputs(4328) <= layer1_outputs(2995);
    layer2_outputs(4329) <= layer1_outputs(1153);
    layer2_outputs(4330) <= layer1_outputs(53);
    layer2_outputs(4331) <= layer1_outputs(9226);
    layer2_outputs(4332) <= not(layer1_outputs(7955)) or (layer1_outputs(5081));
    layer2_outputs(4333) <= not(layer1_outputs(1836));
    layer2_outputs(4334) <= not(layer1_outputs(3340));
    layer2_outputs(4335) <= not(layer1_outputs(3571));
    layer2_outputs(4336) <= not((layer1_outputs(1727)) xor (layer1_outputs(8624)));
    layer2_outputs(4337) <= layer1_outputs(7227);
    layer2_outputs(4338) <= not(layer1_outputs(3953));
    layer2_outputs(4339) <= not(layer1_outputs(9237));
    layer2_outputs(4340) <= not((layer1_outputs(5036)) or (layer1_outputs(4169)));
    layer2_outputs(4341) <= not(layer1_outputs(9213));
    layer2_outputs(4342) <= (layer1_outputs(6118)) and (layer1_outputs(5045));
    layer2_outputs(4343) <= not(layer1_outputs(2920));
    layer2_outputs(4344) <= layer1_outputs(3255);
    layer2_outputs(4345) <= not((layer1_outputs(3332)) or (layer1_outputs(3251)));
    layer2_outputs(4346) <= layer1_outputs(4948);
    layer2_outputs(4347) <= not((layer1_outputs(4891)) xor (layer1_outputs(1834)));
    layer2_outputs(4348) <= not(layer1_outputs(4998));
    layer2_outputs(4349) <= (layer1_outputs(976)) and not (layer1_outputs(869));
    layer2_outputs(4350) <= not(layer1_outputs(5354));
    layer2_outputs(4351) <= not(layer1_outputs(3207));
    layer2_outputs(4352) <= not(layer1_outputs(2717)) or (layer1_outputs(2700));
    layer2_outputs(4353) <= not((layer1_outputs(5046)) xor (layer1_outputs(828)));
    layer2_outputs(4354) <= not((layer1_outputs(1339)) or (layer1_outputs(7395)));
    layer2_outputs(4355) <= (layer1_outputs(8193)) and not (layer1_outputs(2063));
    layer2_outputs(4356) <= not(layer1_outputs(8602)) or (layer1_outputs(9095));
    layer2_outputs(4357) <= layer1_outputs(9675);
    layer2_outputs(4358) <= not((layer1_outputs(10092)) and (layer1_outputs(5591)));
    layer2_outputs(4359) <= not(layer1_outputs(2073));
    layer2_outputs(4360) <= (layer1_outputs(883)) xor (layer1_outputs(2727));
    layer2_outputs(4361) <= not(layer1_outputs(1792));
    layer2_outputs(4362) <= not((layer1_outputs(647)) or (layer1_outputs(6509)));
    layer2_outputs(4363) <= (layer1_outputs(87)) or (layer1_outputs(3193));
    layer2_outputs(4364) <= not(layer1_outputs(3312));
    layer2_outputs(4365) <= layer1_outputs(274);
    layer2_outputs(4366) <= (layer1_outputs(7339)) and not (layer1_outputs(8203));
    layer2_outputs(4367) <= not(layer1_outputs(9387));
    layer2_outputs(4368) <= (layer1_outputs(2998)) and not (layer1_outputs(2865));
    layer2_outputs(4369) <= layer1_outputs(9114);
    layer2_outputs(4370) <= not(layer1_outputs(9014)) or (layer1_outputs(5847));
    layer2_outputs(4371) <= (layer1_outputs(4678)) xor (layer1_outputs(6077));
    layer2_outputs(4372) <= not(layer1_outputs(4337));
    layer2_outputs(4373) <= not(layer1_outputs(4837));
    layer2_outputs(4374) <= (layer1_outputs(6025)) and not (layer1_outputs(9661));
    layer2_outputs(4375) <= not(layer1_outputs(1943));
    layer2_outputs(4376) <= layer1_outputs(9716);
    layer2_outputs(4377) <= layer1_outputs(659);
    layer2_outputs(4378) <= not(layer1_outputs(7951));
    layer2_outputs(4379) <= not(layer1_outputs(2149));
    layer2_outputs(4380) <= (layer1_outputs(840)) xor (layer1_outputs(1081));
    layer2_outputs(4381) <= not(layer1_outputs(2227));
    layer2_outputs(4382) <= layer1_outputs(8357);
    layer2_outputs(4383) <= not(layer1_outputs(6641));
    layer2_outputs(4384) <= not(layer1_outputs(6815)) or (layer1_outputs(4059));
    layer2_outputs(4385) <= (layer1_outputs(5538)) and not (layer1_outputs(3247));
    layer2_outputs(4386) <= layer1_outputs(5085);
    layer2_outputs(4387) <= layer1_outputs(808);
    layer2_outputs(4388) <= layer1_outputs(4348);
    layer2_outputs(4389) <= (layer1_outputs(5225)) and not (layer1_outputs(448));
    layer2_outputs(4390) <= (layer1_outputs(8838)) or (layer1_outputs(6156));
    layer2_outputs(4391) <= (layer1_outputs(3349)) or (layer1_outputs(2875));
    layer2_outputs(4392) <= not(layer1_outputs(934));
    layer2_outputs(4393) <= not((layer1_outputs(1394)) xor (layer1_outputs(1017)));
    layer2_outputs(4394) <= layer1_outputs(4727);
    layer2_outputs(4395) <= layer1_outputs(4841);
    layer2_outputs(4396) <= not(layer1_outputs(2557)) or (layer1_outputs(2131));
    layer2_outputs(4397) <= layer1_outputs(2396);
    layer2_outputs(4398) <= not(layer1_outputs(1024));
    layer2_outputs(4399) <= '1';
    layer2_outputs(4400) <= not(layer1_outputs(5679));
    layer2_outputs(4401) <= (layer1_outputs(1689)) xor (layer1_outputs(2036));
    layer2_outputs(4402) <= layer1_outputs(6432);
    layer2_outputs(4403) <= (layer1_outputs(3093)) and not (layer1_outputs(6893));
    layer2_outputs(4404) <= not((layer1_outputs(3282)) or (layer1_outputs(7837)));
    layer2_outputs(4405) <= not(layer1_outputs(3694)) or (layer1_outputs(8195));
    layer2_outputs(4406) <= (layer1_outputs(6615)) and not (layer1_outputs(3617));
    layer2_outputs(4407) <= (layer1_outputs(5045)) and not (layer1_outputs(9208));
    layer2_outputs(4408) <= not(layer1_outputs(8033)) or (layer1_outputs(9188));
    layer2_outputs(4409) <= not(layer1_outputs(9207));
    layer2_outputs(4410) <= (layer1_outputs(6766)) and not (layer1_outputs(3337));
    layer2_outputs(4411) <= (layer1_outputs(2786)) xor (layer1_outputs(2376));
    layer2_outputs(4412) <= not(layer1_outputs(7889)) or (layer1_outputs(303));
    layer2_outputs(4413) <= layer1_outputs(6312);
    layer2_outputs(4414) <= layer1_outputs(65);
    layer2_outputs(4415) <= not(layer1_outputs(1087));
    layer2_outputs(4416) <= (layer1_outputs(2487)) or (layer1_outputs(6665));
    layer2_outputs(4417) <= not(layer1_outputs(2976));
    layer2_outputs(4418) <= not(layer1_outputs(4398)) or (layer1_outputs(5547));
    layer2_outputs(4419) <= (layer1_outputs(3462)) and not (layer1_outputs(3300));
    layer2_outputs(4420) <= layer1_outputs(2940);
    layer2_outputs(4421) <= (layer1_outputs(9755)) and not (layer1_outputs(8230));
    layer2_outputs(4422) <= (layer1_outputs(415)) or (layer1_outputs(5509));
    layer2_outputs(4423) <= not((layer1_outputs(1386)) or (layer1_outputs(4508)));
    layer2_outputs(4424) <= not(layer1_outputs(2103));
    layer2_outputs(4425) <= not(layer1_outputs(8111));
    layer2_outputs(4426) <= (layer1_outputs(1975)) and not (layer1_outputs(8527));
    layer2_outputs(4427) <= not((layer1_outputs(2323)) or (layer1_outputs(9490)));
    layer2_outputs(4428) <= not((layer1_outputs(8184)) and (layer1_outputs(6082)));
    layer2_outputs(4429) <= '0';
    layer2_outputs(4430) <= not((layer1_outputs(9952)) or (layer1_outputs(7012)));
    layer2_outputs(4431) <= not(layer1_outputs(4752));
    layer2_outputs(4432) <= layer1_outputs(4270);
    layer2_outputs(4433) <= (layer1_outputs(8108)) xor (layer1_outputs(5284));
    layer2_outputs(4434) <= (layer1_outputs(306)) and not (layer1_outputs(1889));
    layer2_outputs(4435) <= (layer1_outputs(7630)) xor (layer1_outputs(69));
    layer2_outputs(4436) <= (layer1_outputs(3069)) and (layer1_outputs(9061));
    layer2_outputs(4437) <= not((layer1_outputs(5194)) xor (layer1_outputs(4250)));
    layer2_outputs(4438) <= (layer1_outputs(1821)) and (layer1_outputs(6304));
    layer2_outputs(4439) <= not((layer1_outputs(4085)) and (layer1_outputs(237)));
    layer2_outputs(4440) <= not((layer1_outputs(2445)) and (layer1_outputs(8359)));
    layer2_outputs(4441) <= layer1_outputs(2061);
    layer2_outputs(4442) <= layer1_outputs(9254);
    layer2_outputs(4443) <= not((layer1_outputs(6343)) or (layer1_outputs(8296)));
    layer2_outputs(4444) <= layer1_outputs(3328);
    layer2_outputs(4445) <= not(layer1_outputs(4178)) or (layer1_outputs(4893));
    layer2_outputs(4446) <= not(layer1_outputs(8145));
    layer2_outputs(4447) <= not((layer1_outputs(1029)) xor (layer1_outputs(4910)));
    layer2_outputs(4448) <= layer1_outputs(5825);
    layer2_outputs(4449) <= layer1_outputs(1001);
    layer2_outputs(4450) <= layer1_outputs(2650);
    layer2_outputs(4451) <= not(layer1_outputs(4049));
    layer2_outputs(4452) <= (layer1_outputs(3917)) and not (layer1_outputs(719));
    layer2_outputs(4453) <= (layer1_outputs(2405)) and not (layer1_outputs(4635));
    layer2_outputs(4454) <= not(layer1_outputs(7116));
    layer2_outputs(4455) <= layer1_outputs(1004);
    layer2_outputs(4456) <= (layer1_outputs(3564)) and not (layer1_outputs(557));
    layer2_outputs(4457) <= (layer1_outputs(1603)) xor (layer1_outputs(3705));
    layer2_outputs(4458) <= not((layer1_outputs(3723)) xor (layer1_outputs(2751)));
    layer2_outputs(4459) <= not(layer1_outputs(5153)) or (layer1_outputs(5090));
    layer2_outputs(4460) <= layer1_outputs(2457);
    layer2_outputs(4461) <= layer1_outputs(9915);
    layer2_outputs(4462) <= not(layer1_outputs(9763));
    layer2_outputs(4463) <= not(layer1_outputs(6409));
    layer2_outputs(4464) <= not((layer1_outputs(7063)) and (layer1_outputs(6817)));
    layer2_outputs(4465) <= not(layer1_outputs(5673));
    layer2_outputs(4466) <= not(layer1_outputs(3418)) or (layer1_outputs(1729));
    layer2_outputs(4467) <= (layer1_outputs(4762)) xor (layer1_outputs(6176));
    layer2_outputs(4468) <= (layer1_outputs(5250)) and not (layer1_outputs(9209));
    layer2_outputs(4469) <= not(layer1_outputs(3863));
    layer2_outputs(4470) <= not(layer1_outputs(2854)) or (layer1_outputs(4168));
    layer2_outputs(4471) <= not((layer1_outputs(1715)) xor (layer1_outputs(1617)));
    layer2_outputs(4472) <= not(layer1_outputs(9783)) or (layer1_outputs(145));
    layer2_outputs(4473) <= layer1_outputs(8640);
    layer2_outputs(4474) <= not(layer1_outputs(6817));
    layer2_outputs(4475) <= layer1_outputs(8254);
    layer2_outputs(4476) <= (layer1_outputs(8725)) and not (layer1_outputs(269));
    layer2_outputs(4477) <= not((layer1_outputs(4330)) and (layer1_outputs(6894)));
    layer2_outputs(4478) <= not((layer1_outputs(7016)) or (layer1_outputs(5180)));
    layer2_outputs(4479) <= not((layer1_outputs(2089)) or (layer1_outputs(13)));
    layer2_outputs(4480) <= layer1_outputs(5144);
    layer2_outputs(4481) <= layer1_outputs(9004);
    layer2_outputs(4482) <= not((layer1_outputs(254)) or (layer1_outputs(10190)));
    layer2_outputs(4483) <= not(layer1_outputs(9101));
    layer2_outputs(4484) <= not(layer1_outputs(6840)) or (layer1_outputs(6758));
    layer2_outputs(4485) <= layer1_outputs(1462);
    layer2_outputs(4486) <= layer1_outputs(10150);
    layer2_outputs(4487) <= layer1_outputs(2862);
    layer2_outputs(4488) <= not(layer1_outputs(5717));
    layer2_outputs(4489) <= not((layer1_outputs(3786)) and (layer1_outputs(8610)));
    layer2_outputs(4490) <= (layer1_outputs(3943)) and (layer1_outputs(8716));
    layer2_outputs(4491) <= layer1_outputs(10122);
    layer2_outputs(4492) <= not(layer1_outputs(4682));
    layer2_outputs(4493) <= not(layer1_outputs(9647));
    layer2_outputs(4494) <= not((layer1_outputs(8447)) or (layer1_outputs(1607)));
    layer2_outputs(4495) <= not(layer1_outputs(5382));
    layer2_outputs(4496) <= not(layer1_outputs(8318));
    layer2_outputs(4497) <= layer1_outputs(1859);
    layer2_outputs(4498) <= '1';
    layer2_outputs(4499) <= layer1_outputs(3447);
    layer2_outputs(4500) <= not((layer1_outputs(6518)) or (layer1_outputs(1076)));
    layer2_outputs(4501) <= not((layer1_outputs(8286)) and (layer1_outputs(6348)));
    layer2_outputs(4502) <= layer1_outputs(6030);
    layer2_outputs(4503) <= layer1_outputs(7828);
    layer2_outputs(4504) <= (layer1_outputs(1989)) and (layer1_outputs(7511));
    layer2_outputs(4505) <= layer1_outputs(1682);
    layer2_outputs(4506) <= (layer1_outputs(73)) xor (layer1_outputs(9064));
    layer2_outputs(4507) <= (layer1_outputs(4179)) and not (layer1_outputs(7613));
    layer2_outputs(4508) <= (layer1_outputs(10126)) and (layer1_outputs(2090));
    layer2_outputs(4509) <= (layer1_outputs(9018)) xor (layer1_outputs(3600));
    layer2_outputs(4510) <= (layer1_outputs(2514)) and not (layer1_outputs(1618));
    layer2_outputs(4511) <= not((layer1_outputs(7104)) and (layer1_outputs(2696)));
    layer2_outputs(4512) <= not(layer1_outputs(1293)) or (layer1_outputs(5572));
    layer2_outputs(4513) <= not(layer1_outputs(4151)) or (layer1_outputs(8294));
    layer2_outputs(4514) <= (layer1_outputs(3246)) xor (layer1_outputs(5975));
    layer2_outputs(4515) <= layer1_outputs(9460);
    layer2_outputs(4516) <= (layer1_outputs(6505)) and (layer1_outputs(5222));
    layer2_outputs(4517) <= layer1_outputs(6613);
    layer2_outputs(4518) <= not(layer1_outputs(3311));
    layer2_outputs(4519) <= (layer1_outputs(8535)) and (layer1_outputs(2759));
    layer2_outputs(4520) <= layer1_outputs(7248);
    layer2_outputs(4521) <= (layer1_outputs(8269)) and (layer1_outputs(6340));
    layer2_outputs(4522) <= layer1_outputs(6704);
    layer2_outputs(4523) <= (layer1_outputs(3727)) and not (layer1_outputs(2292));
    layer2_outputs(4524) <= not(layer1_outputs(7244));
    layer2_outputs(4525) <= not((layer1_outputs(7078)) or (layer1_outputs(6576)));
    layer2_outputs(4526) <= not((layer1_outputs(7967)) xor (layer1_outputs(5829)));
    layer2_outputs(4527) <= (layer1_outputs(5034)) and not (layer1_outputs(6424));
    layer2_outputs(4528) <= (layer1_outputs(4532)) and (layer1_outputs(4602));
    layer2_outputs(4529) <= not(layer1_outputs(8240));
    layer2_outputs(4530) <= layer1_outputs(8069);
    layer2_outputs(4531) <= layer1_outputs(123);
    layer2_outputs(4532) <= not((layer1_outputs(7060)) xor (layer1_outputs(4437)));
    layer2_outputs(4533) <= not(layer1_outputs(1894));
    layer2_outputs(4534) <= not((layer1_outputs(7853)) and (layer1_outputs(3414)));
    layer2_outputs(4535) <= (layer1_outputs(3595)) xor (layer1_outputs(3160));
    layer2_outputs(4536) <= (layer1_outputs(8779)) and (layer1_outputs(7724));
    layer2_outputs(4537) <= layer1_outputs(10117);
    layer2_outputs(4538) <= layer1_outputs(8532);
    layer2_outputs(4539) <= not(layer1_outputs(2770));
    layer2_outputs(4540) <= (layer1_outputs(4499)) and not (layer1_outputs(7099));
    layer2_outputs(4541) <= (layer1_outputs(4013)) and (layer1_outputs(2888));
    layer2_outputs(4542) <= layer1_outputs(458);
    layer2_outputs(4543) <= not(layer1_outputs(1191));
    layer2_outputs(4544) <= not((layer1_outputs(2161)) and (layer1_outputs(3743)));
    layer2_outputs(4545) <= (layer1_outputs(8779)) and (layer1_outputs(1585));
    layer2_outputs(4546) <= not(layer1_outputs(3226)) or (layer1_outputs(7978));
    layer2_outputs(4547) <= not((layer1_outputs(4708)) and (layer1_outputs(3191)));
    layer2_outputs(4548) <= layer1_outputs(9859);
    layer2_outputs(4549) <= (layer1_outputs(6090)) and not (layer1_outputs(5243));
    layer2_outputs(4550) <= layer1_outputs(551);
    layer2_outputs(4551) <= not(layer1_outputs(2124));
    layer2_outputs(4552) <= not(layer1_outputs(5707));
    layer2_outputs(4553) <= layer1_outputs(8243);
    layer2_outputs(4554) <= not(layer1_outputs(5438));
    layer2_outputs(4555) <= not(layer1_outputs(8191)) or (layer1_outputs(10049));
    layer2_outputs(4556) <= layer1_outputs(1559);
    layer2_outputs(4557) <= not((layer1_outputs(3330)) xor (layer1_outputs(10009)));
    layer2_outputs(4558) <= not(layer1_outputs(2455));
    layer2_outputs(4559) <= (layer1_outputs(2104)) and not (layer1_outputs(6606));
    layer2_outputs(4560) <= not(layer1_outputs(503)) or (layer1_outputs(5627));
    layer2_outputs(4561) <= not(layer1_outputs(2220));
    layer2_outputs(4562) <= not(layer1_outputs(1909)) or (layer1_outputs(3151));
    layer2_outputs(4563) <= not((layer1_outputs(116)) xor (layer1_outputs(548)));
    layer2_outputs(4564) <= not(layer1_outputs(2754));
    layer2_outputs(4565) <= not(layer1_outputs(9097));
    layer2_outputs(4566) <= not(layer1_outputs(3033));
    layer2_outputs(4567) <= not((layer1_outputs(1305)) xor (layer1_outputs(5318)));
    layer2_outputs(4568) <= (layer1_outputs(9164)) xor (layer1_outputs(9947));
    layer2_outputs(4569) <= '1';
    layer2_outputs(4570) <= (layer1_outputs(4299)) and (layer1_outputs(7895));
    layer2_outputs(4571) <= layer1_outputs(1937);
    layer2_outputs(4572) <= not((layer1_outputs(1403)) and (layer1_outputs(1132)));
    layer2_outputs(4573) <= layer1_outputs(1758);
    layer2_outputs(4574) <= layer1_outputs(9854);
    layer2_outputs(4575) <= (layer1_outputs(8481)) xor (layer1_outputs(4181));
    layer2_outputs(4576) <= (layer1_outputs(8741)) xor (layer1_outputs(1510));
    layer2_outputs(4577) <= layer1_outputs(870);
    layer2_outputs(4578) <= not((layer1_outputs(9110)) and (layer1_outputs(5052)));
    layer2_outputs(4579) <= layer1_outputs(2102);
    layer2_outputs(4580) <= not(layer1_outputs(6457));
    layer2_outputs(4581) <= not((layer1_outputs(1012)) and (layer1_outputs(4955)));
    layer2_outputs(4582) <= layer1_outputs(8344);
    layer2_outputs(4583) <= not((layer1_outputs(8929)) xor (layer1_outputs(6150)));
    layer2_outputs(4584) <= not(layer1_outputs(4763)) or (layer1_outputs(958));
    layer2_outputs(4585) <= (layer1_outputs(5583)) or (layer1_outputs(2058));
    layer2_outputs(4586) <= (layer1_outputs(7863)) and not (layer1_outputs(8781));
    layer2_outputs(4587) <= not(layer1_outputs(7968));
    layer2_outputs(4588) <= not(layer1_outputs(2665)) or (layer1_outputs(6517));
    layer2_outputs(4589) <= (layer1_outputs(2151)) or (layer1_outputs(2742));
    layer2_outputs(4590) <= (layer1_outputs(1320)) xor (layer1_outputs(1860));
    layer2_outputs(4591) <= not(layer1_outputs(23)) or (layer1_outputs(3211));
    layer2_outputs(4592) <= not((layer1_outputs(6334)) or (layer1_outputs(809)));
    layer2_outputs(4593) <= (layer1_outputs(794)) and not (layer1_outputs(1311));
    layer2_outputs(4594) <= layer1_outputs(3040);
    layer2_outputs(4595) <= (layer1_outputs(3713)) and not (layer1_outputs(8380));
    layer2_outputs(4596) <= not((layer1_outputs(7821)) or (layer1_outputs(6700)));
    layer2_outputs(4597) <= not(layer1_outputs(9364));
    layer2_outputs(4598) <= layer1_outputs(8632);
    layer2_outputs(4599) <= not(layer1_outputs(4282));
    layer2_outputs(4600) <= (layer1_outputs(5796)) and (layer1_outputs(5633));
    layer2_outputs(4601) <= (layer1_outputs(3266)) or (layer1_outputs(52));
    layer2_outputs(4602) <= layer1_outputs(6792);
    layer2_outputs(4603) <= not(layer1_outputs(8598));
    layer2_outputs(4604) <= not((layer1_outputs(1902)) xor (layer1_outputs(655)));
    layer2_outputs(4605) <= not((layer1_outputs(4081)) or (layer1_outputs(5588)));
    layer2_outputs(4606) <= (layer1_outputs(6515)) or (layer1_outputs(8103));
    layer2_outputs(4607) <= layer1_outputs(551);
    layer2_outputs(4608) <= (layer1_outputs(8732)) or (layer1_outputs(2729));
    layer2_outputs(4609) <= not(layer1_outputs(8879));
    layer2_outputs(4610) <= not(layer1_outputs(3764));
    layer2_outputs(4611) <= not((layer1_outputs(543)) xor (layer1_outputs(586)));
    layer2_outputs(4612) <= (layer1_outputs(6028)) and not (layer1_outputs(3531));
    layer2_outputs(4613) <= layer1_outputs(1265);
    layer2_outputs(4614) <= (layer1_outputs(6932)) and not (layer1_outputs(8342));
    layer2_outputs(4615) <= layer1_outputs(1718);
    layer2_outputs(4616) <= layer1_outputs(2092);
    layer2_outputs(4617) <= layer1_outputs(7566);
    layer2_outputs(4618) <= layer1_outputs(2224);
    layer2_outputs(4619) <= not((layer1_outputs(2272)) or (layer1_outputs(2394)));
    layer2_outputs(4620) <= not(layer1_outputs(5742));
    layer2_outputs(4621) <= not((layer1_outputs(2727)) and (layer1_outputs(9920)));
    layer2_outputs(4622) <= layer1_outputs(4340);
    layer2_outputs(4623) <= not((layer1_outputs(3772)) and (layer1_outputs(9089)));
    layer2_outputs(4624) <= not(layer1_outputs(732));
    layer2_outputs(4625) <= (layer1_outputs(1193)) and not (layer1_outputs(641));
    layer2_outputs(4626) <= not((layer1_outputs(10206)) and (layer1_outputs(3336)));
    layer2_outputs(4627) <= not(layer1_outputs(3642)) or (layer1_outputs(7007));
    layer2_outputs(4628) <= not(layer1_outputs(4110));
    layer2_outputs(4629) <= not((layer1_outputs(2545)) xor (layer1_outputs(5705)));
    layer2_outputs(4630) <= not((layer1_outputs(1496)) xor (layer1_outputs(44)));
    layer2_outputs(4631) <= not((layer1_outputs(4637)) or (layer1_outputs(11)));
    layer2_outputs(4632) <= layer1_outputs(2468);
    layer2_outputs(4633) <= layer1_outputs(662);
    layer2_outputs(4634) <= layer1_outputs(5990);
    layer2_outputs(4635) <= layer1_outputs(6165);
    layer2_outputs(4636) <= not(layer1_outputs(5959));
    layer2_outputs(4637) <= not(layer1_outputs(1760));
    layer2_outputs(4638) <= layer1_outputs(6109);
    layer2_outputs(4639) <= not((layer1_outputs(4137)) xor (layer1_outputs(8370)));
    layer2_outputs(4640) <= '0';
    layer2_outputs(4641) <= layer1_outputs(1883);
    layer2_outputs(4642) <= layer1_outputs(9942);
    layer2_outputs(4643) <= not((layer1_outputs(1510)) and (layer1_outputs(7299)));
    layer2_outputs(4644) <= layer1_outputs(7750);
    layer2_outputs(4645) <= (layer1_outputs(2796)) and not (layer1_outputs(4586));
    layer2_outputs(4646) <= layer1_outputs(10226);
    layer2_outputs(4647) <= not(layer1_outputs(4335));
    layer2_outputs(4648) <= not(layer1_outputs(2218));
    layer2_outputs(4649) <= layer1_outputs(3111);
    layer2_outputs(4650) <= not((layer1_outputs(10221)) and (layer1_outputs(3284)));
    layer2_outputs(4651) <= (layer1_outputs(7709)) and not (layer1_outputs(8233));
    layer2_outputs(4652) <= (layer1_outputs(2425)) and (layer1_outputs(5556));
    layer2_outputs(4653) <= (layer1_outputs(4405)) or (layer1_outputs(9551));
    layer2_outputs(4654) <= layer1_outputs(2631);
    layer2_outputs(4655) <= '1';
    layer2_outputs(4656) <= not(layer1_outputs(3109)) or (layer1_outputs(4231));
    layer2_outputs(4657) <= not(layer1_outputs(5509)) or (layer1_outputs(6335));
    layer2_outputs(4658) <= not(layer1_outputs(3243));
    layer2_outputs(4659) <= not(layer1_outputs(2821));
    layer2_outputs(4660) <= (layer1_outputs(4496)) xor (layer1_outputs(5428));
    layer2_outputs(4661) <= not(layer1_outputs(9742));
    layer2_outputs(4662) <= (layer1_outputs(4265)) and not (layer1_outputs(8758));
    layer2_outputs(4663) <= not(layer1_outputs(5098));
    layer2_outputs(4664) <= not(layer1_outputs(8172));
    layer2_outputs(4665) <= (layer1_outputs(8207)) and not (layer1_outputs(7388));
    layer2_outputs(4666) <= layer1_outputs(1298);
    layer2_outputs(4667) <= layer1_outputs(10173);
    layer2_outputs(4668) <= (layer1_outputs(1034)) and (layer1_outputs(6851));
    layer2_outputs(4669) <= layer1_outputs(1588);
    layer2_outputs(4670) <= (layer1_outputs(5340)) and not (layer1_outputs(588));
    layer2_outputs(4671) <= (layer1_outputs(7390)) and (layer1_outputs(3362));
    layer2_outputs(4672) <= not(layer1_outputs(9240)) or (layer1_outputs(7083));
    layer2_outputs(4673) <= layer1_outputs(5151);
    layer2_outputs(4674) <= not(layer1_outputs(7902)) or (layer1_outputs(2300));
    layer2_outputs(4675) <= not(layer1_outputs(3600));
    layer2_outputs(4676) <= layer1_outputs(2469);
    layer2_outputs(4677) <= not(layer1_outputs(3161)) or (layer1_outputs(3454));
    layer2_outputs(4678) <= (layer1_outputs(9791)) xor (layer1_outputs(9580));
    layer2_outputs(4679) <= (layer1_outputs(2266)) xor (layer1_outputs(8017));
    layer2_outputs(4680) <= not(layer1_outputs(4496)) or (layer1_outputs(3135));
    layer2_outputs(4681) <= (layer1_outputs(7467)) xor (layer1_outputs(7321));
    layer2_outputs(4682) <= not(layer1_outputs(1873));
    layer2_outputs(4683) <= layer1_outputs(1379);
    layer2_outputs(4684) <= not(layer1_outputs(5643));
    layer2_outputs(4685) <= not(layer1_outputs(6388));
    layer2_outputs(4686) <= layer1_outputs(5505);
    layer2_outputs(4687) <= (layer1_outputs(4681)) or (layer1_outputs(7146));
    layer2_outputs(4688) <= layer1_outputs(8682);
    layer2_outputs(4689) <= (layer1_outputs(1314)) and not (layer1_outputs(3484));
    layer2_outputs(4690) <= not((layer1_outputs(3581)) xor (layer1_outputs(4453)));
    layer2_outputs(4691) <= not(layer1_outputs(3591)) or (layer1_outputs(6072));
    layer2_outputs(4692) <= (layer1_outputs(8950)) or (layer1_outputs(2789));
    layer2_outputs(4693) <= (layer1_outputs(3232)) and (layer1_outputs(1497));
    layer2_outputs(4694) <= not(layer1_outputs(6348)) or (layer1_outputs(3741));
    layer2_outputs(4695) <= (layer1_outputs(7657)) and not (layer1_outputs(789));
    layer2_outputs(4696) <= not(layer1_outputs(1681));
    layer2_outputs(4697) <= (layer1_outputs(3399)) and not (layer1_outputs(6055));
    layer2_outputs(4698) <= (layer1_outputs(642)) and not (layer1_outputs(365));
    layer2_outputs(4699) <= not(layer1_outputs(9470));
    layer2_outputs(4700) <= not(layer1_outputs(7255)) or (layer1_outputs(2656));
    layer2_outputs(4701) <= (layer1_outputs(5275)) xor (layer1_outputs(3618));
    layer2_outputs(4702) <= not(layer1_outputs(4673));
    layer2_outputs(4703) <= layer1_outputs(9770);
    layer2_outputs(4704) <= not(layer1_outputs(5901));
    layer2_outputs(4705) <= layer1_outputs(6429);
    layer2_outputs(4706) <= not(layer1_outputs(4970));
    layer2_outputs(4707) <= layer1_outputs(4402);
    layer2_outputs(4708) <= (layer1_outputs(4739)) or (layer1_outputs(5590));
    layer2_outputs(4709) <= layer1_outputs(1855);
    layer2_outputs(4710) <= not(layer1_outputs(1269)) or (layer1_outputs(2598));
    layer2_outputs(4711) <= not((layer1_outputs(3355)) or (layer1_outputs(6262)));
    layer2_outputs(4712) <= layer1_outputs(718);
    layer2_outputs(4713) <= not(layer1_outputs(3029));
    layer2_outputs(4714) <= (layer1_outputs(3007)) and (layer1_outputs(3691));
    layer2_outputs(4715) <= not(layer1_outputs(275)) or (layer1_outputs(4943));
    layer2_outputs(4716) <= not(layer1_outputs(2214)) or (layer1_outputs(9787));
    layer2_outputs(4717) <= not((layer1_outputs(1803)) and (layer1_outputs(7857)));
    layer2_outputs(4718) <= not(layer1_outputs(3601));
    layer2_outputs(4719) <= layer1_outputs(981);
    layer2_outputs(4720) <= layer1_outputs(4212);
    layer2_outputs(4721) <= (layer1_outputs(8572)) and (layer1_outputs(1349));
    layer2_outputs(4722) <= not(layer1_outputs(6308));
    layer2_outputs(4723) <= not((layer1_outputs(3099)) or (layer1_outputs(5566)));
    layer2_outputs(4724) <= (layer1_outputs(1900)) xor (layer1_outputs(369));
    layer2_outputs(4725) <= (layer1_outputs(783)) and (layer1_outputs(2698));
    layer2_outputs(4726) <= not(layer1_outputs(879));
    layer2_outputs(4727) <= not(layer1_outputs(1451));
    layer2_outputs(4728) <= layer1_outputs(3309);
    layer2_outputs(4729) <= (layer1_outputs(8365)) and not (layer1_outputs(5639));
    layer2_outputs(4730) <= (layer1_outputs(9383)) and (layer1_outputs(3783));
    layer2_outputs(4731) <= layer1_outputs(9696);
    layer2_outputs(4732) <= not((layer1_outputs(2725)) xor (layer1_outputs(4933)));
    layer2_outputs(4733) <= not(layer1_outputs(32));
    layer2_outputs(4734) <= (layer1_outputs(8293)) xor (layer1_outputs(1893));
    layer2_outputs(4735) <= (layer1_outputs(9662)) xor (layer1_outputs(8773));
    layer2_outputs(4736) <= not(layer1_outputs(6446)) or (layer1_outputs(5393));
    layer2_outputs(4737) <= not(layer1_outputs(6112)) or (layer1_outputs(8153));
    layer2_outputs(4738) <= not((layer1_outputs(590)) xor (layer1_outputs(6127)));
    layer2_outputs(4739) <= not(layer1_outputs(3824));
    layer2_outputs(4740) <= layer1_outputs(1353);
    layer2_outputs(4741) <= not((layer1_outputs(4246)) xor (layer1_outputs(9798)));
    layer2_outputs(4742) <= not(layer1_outputs(7908));
    layer2_outputs(4743) <= not(layer1_outputs(9702));
    layer2_outputs(4744) <= not((layer1_outputs(5471)) or (layer1_outputs(7337)));
    layer2_outputs(4745) <= not((layer1_outputs(4254)) or (layer1_outputs(4288)));
    layer2_outputs(4746) <= layer1_outputs(895);
    layer2_outputs(4747) <= layer1_outputs(1455);
    layer2_outputs(4748) <= (layer1_outputs(1294)) and (layer1_outputs(1052));
    layer2_outputs(4749) <= not(layer1_outputs(1896));
    layer2_outputs(4750) <= not((layer1_outputs(2067)) and (layer1_outputs(2893)));
    layer2_outputs(4751) <= layer1_outputs(7703);
    layer2_outputs(4752) <= layer1_outputs(3730);
    layer2_outputs(4753) <= not(layer1_outputs(429));
    layer2_outputs(4754) <= not((layer1_outputs(6682)) xor (layer1_outputs(4314)));
    layer2_outputs(4755) <= layer1_outputs(4218);
    layer2_outputs(4756) <= (layer1_outputs(8005)) and not (layer1_outputs(764));
    layer2_outputs(4757) <= not((layer1_outputs(3971)) or (layer1_outputs(4281)));
    layer2_outputs(4758) <= layer1_outputs(7951);
    layer2_outputs(4759) <= layer1_outputs(1374);
    layer2_outputs(4760) <= layer1_outputs(1236);
    layer2_outputs(4761) <= not((layer1_outputs(8164)) xor (layer1_outputs(1368)));
    layer2_outputs(4762) <= layer1_outputs(4381);
    layer2_outputs(4763) <= not(layer1_outputs(867));
    layer2_outputs(4764) <= layer1_outputs(2648);
    layer2_outputs(4765) <= layer1_outputs(7383);
    layer2_outputs(4766) <= (layer1_outputs(4688)) or (layer1_outputs(3925));
    layer2_outputs(4767) <= layer1_outputs(5869);
    layer2_outputs(4768) <= not(layer1_outputs(36)) or (layer1_outputs(3488));
    layer2_outputs(4769) <= not(layer1_outputs(5000));
    layer2_outputs(4770) <= (layer1_outputs(157)) or (layer1_outputs(3622));
    layer2_outputs(4771) <= not(layer1_outputs(877));
    layer2_outputs(4772) <= not(layer1_outputs(729));
    layer2_outputs(4773) <= not(layer1_outputs(1084));
    layer2_outputs(4774) <= layer1_outputs(4298);
    layer2_outputs(4775) <= (layer1_outputs(1125)) or (layer1_outputs(9742));
    layer2_outputs(4776) <= not((layer1_outputs(7757)) xor (layer1_outputs(4271)));
    layer2_outputs(4777) <= (layer1_outputs(6647)) xor (layer1_outputs(1036));
    layer2_outputs(4778) <= (layer1_outputs(1389)) or (layer1_outputs(7512));
    layer2_outputs(4779) <= (layer1_outputs(7380)) and not (layer1_outputs(9141));
    layer2_outputs(4780) <= not(layer1_outputs(9164));
    layer2_outputs(4781) <= not(layer1_outputs(8384));
    layer2_outputs(4782) <= not(layer1_outputs(7613));
    layer2_outputs(4783) <= not(layer1_outputs(291));
    layer2_outputs(4784) <= layer1_outputs(6012);
    layer2_outputs(4785) <= not(layer1_outputs(10080));
    layer2_outputs(4786) <= not(layer1_outputs(10145)) or (layer1_outputs(6522));
    layer2_outputs(4787) <= not(layer1_outputs(2105));
    layer2_outputs(4788) <= (layer1_outputs(2637)) or (layer1_outputs(6461));
    layer2_outputs(4789) <= (layer1_outputs(8553)) or (layer1_outputs(2382));
    layer2_outputs(4790) <= not(layer1_outputs(523));
    layer2_outputs(4791) <= (layer1_outputs(9981)) and (layer1_outputs(1776));
    layer2_outputs(4792) <= not((layer1_outputs(3013)) or (layer1_outputs(7173)));
    layer2_outputs(4793) <= not((layer1_outputs(5949)) xor (layer1_outputs(10171)));
    layer2_outputs(4794) <= not(layer1_outputs(5800));
    layer2_outputs(4795) <= (layer1_outputs(5662)) or (layer1_outputs(652));
    layer2_outputs(4796) <= not(layer1_outputs(2807));
    layer2_outputs(4797) <= (layer1_outputs(2349)) and not (layer1_outputs(4725));
    layer2_outputs(4798) <= layer1_outputs(1703);
    layer2_outputs(4799) <= not(layer1_outputs(8104)) or (layer1_outputs(6224));
    layer2_outputs(4800) <= (layer1_outputs(4131)) xor (layer1_outputs(4745));
    layer2_outputs(4801) <= not((layer1_outputs(9298)) and (layer1_outputs(8469)));
    layer2_outputs(4802) <= (layer1_outputs(1240)) and not (layer1_outputs(8476));
    layer2_outputs(4803) <= not(layer1_outputs(9917));
    layer2_outputs(4804) <= (layer1_outputs(8594)) and not (layer1_outputs(5160));
    layer2_outputs(4805) <= layer1_outputs(3252);
    layer2_outputs(4806) <= (layer1_outputs(6373)) and not (layer1_outputs(632));
    layer2_outputs(4807) <= layer1_outputs(1629);
    layer2_outputs(4808) <= not((layer1_outputs(2860)) and (layer1_outputs(1800)));
    layer2_outputs(4809) <= layer1_outputs(9835);
    layer2_outputs(4810) <= not(layer1_outputs(7852)) or (layer1_outputs(4119));
    layer2_outputs(4811) <= layer1_outputs(4389);
    layer2_outputs(4812) <= not(layer1_outputs(8329));
    layer2_outputs(4813) <= not((layer1_outputs(4974)) or (layer1_outputs(5652)));
    layer2_outputs(4814) <= not(layer1_outputs(1228)) or (layer1_outputs(240));
    layer2_outputs(4815) <= not(layer1_outputs(7216));
    layer2_outputs(4816) <= layer1_outputs(433);
    layer2_outputs(4817) <= '1';
    layer2_outputs(4818) <= not(layer1_outputs(3333));
    layer2_outputs(4819) <= not(layer1_outputs(6610)) or (layer1_outputs(9077));
    layer2_outputs(4820) <= not(layer1_outputs(9180)) or (layer1_outputs(1613));
    layer2_outputs(4821) <= layer1_outputs(5771);
    layer2_outputs(4822) <= not(layer1_outputs(9209)) or (layer1_outputs(4698));
    layer2_outputs(4823) <= (layer1_outputs(279)) and not (layer1_outputs(2268));
    layer2_outputs(4824) <= (layer1_outputs(2657)) or (layer1_outputs(9697));
    layer2_outputs(4825) <= not(layer1_outputs(8733)) or (layer1_outputs(5899));
    layer2_outputs(4826) <= not(layer1_outputs(6391));
    layer2_outputs(4827) <= (layer1_outputs(3062)) and not (layer1_outputs(5592));
    layer2_outputs(4828) <= layer1_outputs(6052);
    layer2_outputs(4829) <= not((layer1_outputs(4554)) and (layer1_outputs(7439)));
    layer2_outputs(4830) <= (layer1_outputs(3823)) and (layer1_outputs(495));
    layer2_outputs(4831) <= not(layer1_outputs(7621));
    layer2_outputs(4832) <= layer1_outputs(4044);
    layer2_outputs(4833) <= (layer1_outputs(838)) and not (layer1_outputs(8665));
    layer2_outputs(4834) <= not(layer1_outputs(7722));
    layer2_outputs(4835) <= not(layer1_outputs(6684));
    layer2_outputs(4836) <= not(layer1_outputs(2059));
    layer2_outputs(4837) <= not((layer1_outputs(8410)) and (layer1_outputs(4883)));
    layer2_outputs(4838) <= layer1_outputs(3855);
    layer2_outputs(4839) <= not((layer1_outputs(10069)) and (layer1_outputs(3087)));
    layer2_outputs(4840) <= layer1_outputs(2724);
    layer2_outputs(4841) <= not((layer1_outputs(1998)) or (layer1_outputs(4934)));
    layer2_outputs(4842) <= not(layer1_outputs(952)) or (layer1_outputs(4464));
    layer2_outputs(4843) <= not(layer1_outputs(10144));
    layer2_outputs(4844) <= (layer1_outputs(8633)) or (layer1_outputs(6718));
    layer2_outputs(4845) <= layer1_outputs(6847);
    layer2_outputs(4846) <= not(layer1_outputs(3016));
    layer2_outputs(4847) <= layer1_outputs(2105);
    layer2_outputs(4848) <= not(layer1_outputs(38));
    layer2_outputs(4849) <= not((layer1_outputs(9246)) or (layer1_outputs(5555)));
    layer2_outputs(4850) <= layer1_outputs(4718);
    layer2_outputs(4851) <= layer1_outputs(448);
    layer2_outputs(4852) <= layer1_outputs(1989);
    layer2_outputs(4853) <= (layer1_outputs(3030)) or (layer1_outputs(7364));
    layer2_outputs(4854) <= layer1_outputs(985);
    layer2_outputs(4855) <= layer1_outputs(4937);
    layer2_outputs(4856) <= not(layer1_outputs(9888));
    layer2_outputs(4857) <= not(layer1_outputs(52)) or (layer1_outputs(1411));
    layer2_outputs(4858) <= (layer1_outputs(1264)) and not (layer1_outputs(2342));
    layer2_outputs(4859) <= not(layer1_outputs(364));
    layer2_outputs(4860) <= not(layer1_outputs(1882));
    layer2_outputs(4861) <= not((layer1_outputs(4774)) xor (layer1_outputs(9281)));
    layer2_outputs(4862) <= not((layer1_outputs(7431)) or (layer1_outputs(6145)));
    layer2_outputs(4863) <= (layer1_outputs(1025)) and not (layer1_outputs(5631));
    layer2_outputs(4864) <= not(layer1_outputs(1105));
    layer2_outputs(4865) <= not((layer1_outputs(3206)) and (layer1_outputs(2579)));
    layer2_outputs(4866) <= (layer1_outputs(1144)) and (layer1_outputs(5080));
    layer2_outputs(4867) <= not(layer1_outputs(249));
    layer2_outputs(4868) <= (layer1_outputs(2573)) and not (layer1_outputs(4497));
    layer2_outputs(4869) <= not((layer1_outputs(9389)) and (layer1_outputs(4197)));
    layer2_outputs(4870) <= not((layer1_outputs(2126)) or (layer1_outputs(3244)));
    layer2_outputs(4871) <= (layer1_outputs(5768)) and (layer1_outputs(2568));
    layer2_outputs(4872) <= layer1_outputs(2833);
    layer2_outputs(4873) <= not(layer1_outputs(2307)) or (layer1_outputs(6842));
    layer2_outputs(4874) <= layer1_outputs(8710);
    layer2_outputs(4875) <= (layer1_outputs(3954)) or (layer1_outputs(4092));
    layer2_outputs(4876) <= not(layer1_outputs(1592));
    layer2_outputs(4877) <= layer1_outputs(6078);
    layer2_outputs(4878) <= not(layer1_outputs(786)) or (layer1_outputs(2580));
    layer2_outputs(4879) <= not(layer1_outputs(6226));
    layer2_outputs(4880) <= not(layer1_outputs(920));
    layer2_outputs(4881) <= (layer1_outputs(618)) and not (layer1_outputs(5088));
    layer2_outputs(4882) <= not((layer1_outputs(3572)) and (layer1_outputs(7213)));
    layer2_outputs(4883) <= not((layer1_outputs(7030)) xor (layer1_outputs(780)));
    layer2_outputs(4884) <= (layer1_outputs(4506)) and not (layer1_outputs(2973));
    layer2_outputs(4885) <= not(layer1_outputs(2190));
    layer2_outputs(4886) <= layer1_outputs(4209);
    layer2_outputs(4887) <= not(layer1_outputs(2255));
    layer2_outputs(4888) <= (layer1_outputs(7357)) or (layer1_outputs(6779));
    layer2_outputs(4889) <= layer1_outputs(3272);
    layer2_outputs(4890) <= not((layer1_outputs(990)) and (layer1_outputs(2501)));
    layer2_outputs(4891) <= (layer1_outputs(2751)) and not (layer1_outputs(281));
    layer2_outputs(4892) <= not(layer1_outputs(5943));
    layer2_outputs(4893) <= (layer1_outputs(2391)) and (layer1_outputs(668));
    layer2_outputs(4894) <= not((layer1_outputs(673)) xor (layer1_outputs(1321)));
    layer2_outputs(4895) <= not((layer1_outputs(6304)) xor (layer1_outputs(7585)));
    layer2_outputs(4896) <= layer1_outputs(4601);
    layer2_outputs(4897) <= layer1_outputs(3129);
    layer2_outputs(4898) <= layer1_outputs(2551);
    layer2_outputs(4899) <= not(layer1_outputs(7929)) or (layer1_outputs(9021));
    layer2_outputs(4900) <= (layer1_outputs(3094)) or (layer1_outputs(243));
    layer2_outputs(4901) <= (layer1_outputs(6466)) and not (layer1_outputs(6463));
    layer2_outputs(4902) <= not(layer1_outputs(1423));
    layer2_outputs(4903) <= not(layer1_outputs(6504));
    layer2_outputs(4904) <= not((layer1_outputs(5508)) xor (layer1_outputs(8578)));
    layer2_outputs(4905) <= layer1_outputs(6838);
    layer2_outputs(4906) <= layer1_outputs(4553);
    layer2_outputs(4907) <= not(layer1_outputs(9792)) or (layer1_outputs(2316));
    layer2_outputs(4908) <= (layer1_outputs(7416)) and not (layer1_outputs(5821));
    layer2_outputs(4909) <= not(layer1_outputs(9975)) or (layer1_outputs(6022));
    layer2_outputs(4910) <= not((layer1_outputs(1851)) or (layer1_outputs(3785)));
    layer2_outputs(4911) <= layer1_outputs(3398);
    layer2_outputs(4912) <= (layer1_outputs(1487)) or (layer1_outputs(471));
    layer2_outputs(4913) <= layer1_outputs(6007);
    layer2_outputs(4914) <= layer1_outputs(1166);
    layer2_outputs(4915) <= not(layer1_outputs(5335)) or (layer1_outputs(7250));
    layer2_outputs(4916) <= (layer1_outputs(5169)) or (layer1_outputs(9811));
    layer2_outputs(4917) <= not((layer1_outputs(848)) or (layer1_outputs(2175)));
    layer2_outputs(4918) <= (layer1_outputs(7751)) and not (layer1_outputs(3889));
    layer2_outputs(4919) <= (layer1_outputs(9396)) or (layer1_outputs(4803));
    layer2_outputs(4920) <= layer1_outputs(6212);
    layer2_outputs(4921) <= layer1_outputs(9455);
    layer2_outputs(4922) <= not(layer1_outputs(9398));
    layer2_outputs(4923) <= not(layer1_outputs(5924));
    layer2_outputs(4924) <= (layer1_outputs(5242)) and (layer1_outputs(8826));
    layer2_outputs(4925) <= layer1_outputs(4724);
    layer2_outputs(4926) <= not((layer1_outputs(7578)) xor (layer1_outputs(5618)));
    layer2_outputs(4927) <= not(layer1_outputs(6760));
    layer2_outputs(4928) <= (layer1_outputs(725)) xor (layer1_outputs(7526));
    layer2_outputs(4929) <= not(layer1_outputs(5262));
    layer2_outputs(4930) <= (layer1_outputs(4966)) or (layer1_outputs(1569));
    layer2_outputs(4931) <= layer1_outputs(1758);
    layer2_outputs(4932) <= not(layer1_outputs(7595));
    layer2_outputs(4933) <= not(layer1_outputs(397)) or (layer1_outputs(6745));
    layer2_outputs(4934) <= not((layer1_outputs(6179)) xor (layer1_outputs(6570)));
    layer2_outputs(4935) <= not(layer1_outputs(8667));
    layer2_outputs(4936) <= (layer1_outputs(2216)) xor (layer1_outputs(6407));
    layer2_outputs(4937) <= not(layer1_outputs(7644));
    layer2_outputs(4938) <= layer1_outputs(8643);
    layer2_outputs(4939) <= not((layer1_outputs(7118)) and (layer1_outputs(1799)));
    layer2_outputs(4940) <= layer1_outputs(3845);
    layer2_outputs(4941) <= (layer1_outputs(7310)) and not (layer1_outputs(517));
    layer2_outputs(4942) <= not(layer1_outputs(4664));
    layer2_outputs(4943) <= not(layer1_outputs(8845));
    layer2_outputs(4944) <= layer1_outputs(2512);
    layer2_outputs(4945) <= not(layer1_outputs(505));
    layer2_outputs(4946) <= not(layer1_outputs(6149));
    layer2_outputs(4947) <= layer1_outputs(10147);
    layer2_outputs(4948) <= layer1_outputs(5673);
    layer2_outputs(4949) <= layer1_outputs(1143);
    layer2_outputs(4950) <= layer1_outputs(4645);
    layer2_outputs(4951) <= not(layer1_outputs(6310));
    layer2_outputs(4952) <= layer1_outputs(6068);
    layer2_outputs(4953) <= layer1_outputs(7916);
    layer2_outputs(4954) <= not(layer1_outputs(3686));
    layer2_outputs(4955) <= not((layer1_outputs(5131)) or (layer1_outputs(9311)));
    layer2_outputs(4956) <= (layer1_outputs(6729)) and (layer1_outputs(9663));
    layer2_outputs(4957) <= not((layer1_outputs(5027)) and (layer1_outputs(9628)));
    layer2_outputs(4958) <= not(layer1_outputs(3911));
    layer2_outputs(4959) <= (layer1_outputs(6952)) xor (layer1_outputs(1952));
    layer2_outputs(4960) <= not(layer1_outputs(4261));
    layer2_outputs(4961) <= layer1_outputs(1796);
    layer2_outputs(4962) <= not(layer1_outputs(9430));
    layer2_outputs(4963) <= not(layer1_outputs(3278)) or (layer1_outputs(391));
    layer2_outputs(4964) <= not(layer1_outputs(3283));
    layer2_outputs(4965) <= not(layer1_outputs(2107));
    layer2_outputs(4966) <= layer1_outputs(1722);
    layer2_outputs(4967) <= layer1_outputs(7248);
    layer2_outputs(4968) <= not((layer1_outputs(420)) xor (layer1_outputs(6123)));
    layer2_outputs(4969) <= layer1_outputs(5992);
    layer2_outputs(4970) <= layer1_outputs(6977);
    layer2_outputs(4971) <= not(layer1_outputs(185)) or (layer1_outputs(7681));
    layer2_outputs(4972) <= (layer1_outputs(9721)) and not (layer1_outputs(2320));
    layer2_outputs(4973) <= layer1_outputs(10013);
    layer2_outputs(4974) <= not(layer1_outputs(2325)) or (layer1_outputs(1408));
    layer2_outputs(4975) <= not((layer1_outputs(1202)) xor (layer1_outputs(1922)));
    layer2_outputs(4976) <= not(layer1_outputs(2497));
    layer2_outputs(4977) <= not(layer1_outputs(2978));
    layer2_outputs(4978) <= (layer1_outputs(1491)) and (layer1_outputs(3128));
    layer2_outputs(4979) <= not((layer1_outputs(9984)) or (layer1_outputs(4638)));
    layer2_outputs(4980) <= not(layer1_outputs(1476)) or (layer1_outputs(9013));
    layer2_outputs(4981) <= layer1_outputs(3378);
    layer2_outputs(4982) <= not(layer1_outputs(2486)) or (layer1_outputs(3793));
    layer2_outputs(4983) <= layer1_outputs(5493);
    layer2_outputs(4984) <= (layer1_outputs(406)) or (layer1_outputs(3108));
    layer2_outputs(4985) <= not(layer1_outputs(9667));
    layer2_outputs(4986) <= layer1_outputs(921);
    layer2_outputs(4987) <= layer1_outputs(9934);
    layer2_outputs(4988) <= not(layer1_outputs(9982)) or (layer1_outputs(3715));
    layer2_outputs(4989) <= layer1_outputs(1691);
    layer2_outputs(4990) <= layer1_outputs(3807);
    layer2_outputs(4991) <= not((layer1_outputs(8097)) and (layer1_outputs(10050)));
    layer2_outputs(4992) <= (layer1_outputs(503)) xor (layer1_outputs(1667));
    layer2_outputs(4993) <= (layer1_outputs(6035)) and not (layer1_outputs(8031));
    layer2_outputs(4994) <= not(layer1_outputs(3438));
    layer2_outputs(4995) <= not((layer1_outputs(3562)) and (layer1_outputs(3982)));
    layer2_outputs(4996) <= not(layer1_outputs(6970));
    layer2_outputs(4997) <= layer1_outputs(7333);
    layer2_outputs(4998) <= (layer1_outputs(6514)) and (layer1_outputs(7576));
    layer2_outputs(4999) <= not((layer1_outputs(1505)) or (layer1_outputs(1555)));
    layer2_outputs(5000) <= layer1_outputs(8801);
    layer2_outputs(5001) <= (layer1_outputs(2980)) and not (layer1_outputs(2003));
    layer2_outputs(5002) <= layer1_outputs(8899);
    layer2_outputs(5003) <= layer1_outputs(2991);
    layer2_outputs(5004) <= layer1_outputs(307);
    layer2_outputs(5005) <= not(layer1_outputs(650));
    layer2_outputs(5006) <= layer1_outputs(3142);
    layer2_outputs(5007) <= not(layer1_outputs(8668));
    layer2_outputs(5008) <= layer1_outputs(2014);
    layer2_outputs(5009) <= not((layer1_outputs(4256)) and (layer1_outputs(6030)));
    layer2_outputs(5010) <= layer1_outputs(1570);
    layer2_outputs(5011) <= layer1_outputs(3825);
    layer2_outputs(5012) <= not(layer1_outputs(10022));
    layer2_outputs(5013) <= not(layer1_outputs(1111));
    layer2_outputs(5014) <= not((layer1_outputs(6476)) or (layer1_outputs(3630)));
    layer2_outputs(5015) <= (layer1_outputs(4657)) and (layer1_outputs(1636));
    layer2_outputs(5016) <= (layer1_outputs(4407)) or (layer1_outputs(1183));
    layer2_outputs(5017) <= not((layer1_outputs(1071)) and (layer1_outputs(3613)));
    layer2_outputs(5018) <= not(layer1_outputs(6525));
    layer2_outputs(5019) <= layer1_outputs(3284);
    layer2_outputs(5020) <= not(layer1_outputs(8653));
    layer2_outputs(5021) <= not(layer1_outputs(4482));
    layer2_outputs(5022) <= layer1_outputs(2735);
    layer2_outputs(5023) <= not((layer1_outputs(648)) xor (layer1_outputs(9525)));
    layer2_outputs(5024) <= layer1_outputs(2676);
    layer2_outputs(5025) <= (layer1_outputs(7594)) and not (layer1_outputs(1104));
    layer2_outputs(5026) <= not(layer1_outputs(4726));
    layer2_outputs(5027) <= (layer1_outputs(6579)) and not (layer1_outputs(6046));
    layer2_outputs(5028) <= not((layer1_outputs(9728)) and (layer1_outputs(1526)));
    layer2_outputs(5029) <= (layer1_outputs(4257)) xor (layer1_outputs(7927));
    layer2_outputs(5030) <= (layer1_outputs(1156)) and not (layer1_outputs(5291));
    layer2_outputs(5031) <= (layer1_outputs(7850)) and not (layer1_outputs(7906));
    layer2_outputs(5032) <= not(layer1_outputs(3130)) or (layer1_outputs(7954));
    layer2_outputs(5033) <= (layer1_outputs(4820)) and not (layer1_outputs(3257));
    layer2_outputs(5034) <= not(layer1_outputs(1824)) or (layer1_outputs(10230));
    layer2_outputs(5035) <= layer1_outputs(5736);
    layer2_outputs(5036) <= not(layer1_outputs(2115)) or (layer1_outputs(364));
    layer2_outputs(5037) <= (layer1_outputs(4830)) or (layer1_outputs(9197));
    layer2_outputs(5038) <= (layer1_outputs(6061)) xor (layer1_outputs(7040));
    layer2_outputs(5039) <= not((layer1_outputs(2161)) and (layer1_outputs(7122)));
    layer2_outputs(5040) <= not((layer1_outputs(5167)) xor (layer1_outputs(2144)));
    layer2_outputs(5041) <= not(layer1_outputs(4888)) or (layer1_outputs(9852));
    layer2_outputs(5042) <= layer1_outputs(1826);
    layer2_outputs(5043) <= not(layer1_outputs(4975));
    layer2_outputs(5044) <= '1';
    layer2_outputs(5045) <= not((layer1_outputs(7836)) xor (layer1_outputs(9731)));
    layer2_outputs(5046) <= '1';
    layer2_outputs(5047) <= (layer1_outputs(1694)) and not (layer1_outputs(4484));
    layer2_outputs(5048) <= not((layer1_outputs(8789)) and (layer1_outputs(8815)));
    layer2_outputs(5049) <= not(layer1_outputs(5444));
    layer2_outputs(5050) <= not(layer1_outputs(6180)) or (layer1_outputs(4675));
    layer2_outputs(5051) <= layer1_outputs(4432);
    layer2_outputs(5052) <= not((layer1_outputs(6240)) and (layer1_outputs(2945)));
    layer2_outputs(5053) <= not((layer1_outputs(7545)) xor (layer1_outputs(7247)));
    layer2_outputs(5054) <= not((layer1_outputs(3020)) xor (layer1_outputs(2108)));
    layer2_outputs(5055) <= not(layer1_outputs(666));
    layer2_outputs(5056) <= (layer1_outputs(7689)) or (layer1_outputs(9160));
    layer2_outputs(5057) <= not(layer1_outputs(3077));
    layer2_outputs(5058) <= not(layer1_outputs(3939));
    layer2_outputs(5059) <= not((layer1_outputs(6604)) or (layer1_outputs(1493)));
    layer2_outputs(5060) <= not(layer1_outputs(3809));
    layer2_outputs(5061) <= layer1_outputs(4174);
    layer2_outputs(5062) <= (layer1_outputs(1168)) or (layer1_outputs(6632));
    layer2_outputs(5063) <= not(layer1_outputs(3818));
    layer2_outputs(5064) <= layer1_outputs(1650);
    layer2_outputs(5065) <= not(layer1_outputs(2054)) or (layer1_outputs(3249));
    layer2_outputs(5066) <= (layer1_outputs(5974)) and not (layer1_outputs(2848));
    layer2_outputs(5067) <= not((layer1_outputs(8669)) xor (layer1_outputs(7229)));
    layer2_outputs(5068) <= not(layer1_outputs(3127));
    layer2_outputs(5069) <= (layer1_outputs(6795)) and not (layer1_outputs(8546));
    layer2_outputs(5070) <= not((layer1_outputs(1561)) xor (layer1_outputs(1859)));
    layer2_outputs(5071) <= layer1_outputs(8189);
    layer2_outputs(5072) <= not(layer1_outputs(8545));
    layer2_outputs(5073) <= layer1_outputs(1245);
    layer2_outputs(5074) <= not((layer1_outputs(5493)) and (layer1_outputs(9631)));
    layer2_outputs(5075) <= not(layer1_outputs(10152));
    layer2_outputs(5076) <= not((layer1_outputs(1807)) and (layer1_outputs(1386)));
    layer2_outputs(5077) <= not((layer1_outputs(1617)) xor (layer1_outputs(5111)));
    layer2_outputs(5078) <= layer1_outputs(4914);
    layer2_outputs(5079) <= not(layer1_outputs(3965)) or (layer1_outputs(131));
    layer2_outputs(5080) <= (layer1_outputs(3890)) and not (layer1_outputs(6538));
    layer2_outputs(5081) <= layer1_outputs(3168);
    layer2_outputs(5082) <= (layer1_outputs(3654)) and not (layer1_outputs(4920));
    layer2_outputs(5083) <= not(layer1_outputs(3100)) or (layer1_outputs(9160));
    layer2_outputs(5084) <= not(layer1_outputs(5510));
    layer2_outputs(5085) <= (layer1_outputs(6294)) xor (layer1_outputs(4339));
    layer2_outputs(5086) <= not(layer1_outputs(1137));
    layer2_outputs(5087) <= layer1_outputs(7219);
    layer2_outputs(5088) <= not((layer1_outputs(3132)) xor (layer1_outputs(1370)));
    layer2_outputs(5089) <= layer1_outputs(8222);
    layer2_outputs(5090) <= not(layer1_outputs(8539));
    layer2_outputs(5091) <= layer1_outputs(10113);
    layer2_outputs(5092) <= not((layer1_outputs(1584)) and (layer1_outputs(2567)));
    layer2_outputs(5093) <= not((layer1_outputs(5755)) and (layer1_outputs(8902)));
    layer2_outputs(5094) <= not(layer1_outputs(9666));
    layer2_outputs(5095) <= not(layer1_outputs(1776)) or (layer1_outputs(9081));
    layer2_outputs(5096) <= not(layer1_outputs(3050));
    layer2_outputs(5097) <= not(layer1_outputs(7761));
    layer2_outputs(5098) <= layer1_outputs(7927);
    layer2_outputs(5099) <= not(layer1_outputs(9749)) or (layer1_outputs(7652));
    layer2_outputs(5100) <= (layer1_outputs(3231)) xor (layer1_outputs(3345));
    layer2_outputs(5101) <= layer1_outputs(2761);
    layer2_outputs(5102) <= (layer1_outputs(5029)) and not (layer1_outputs(4926));
    layer2_outputs(5103) <= layer1_outputs(8935);
    layer2_outputs(5104) <= not(layer1_outputs(9150));
    layer2_outputs(5105) <= (layer1_outputs(3682)) and not (layer1_outputs(1740));
    layer2_outputs(5106) <= not(layer1_outputs(7410));
    layer2_outputs(5107) <= layer1_outputs(9980);
    layer2_outputs(5108) <= not(layer1_outputs(5816));
    layer2_outputs(5109) <= layer1_outputs(2482);
    layer2_outputs(5110) <= (layer1_outputs(10041)) xor (layer1_outputs(7694));
    layer2_outputs(5111) <= not(layer1_outputs(3762));
    layer2_outputs(5112) <= (layer1_outputs(1304)) and not (layer1_outputs(5270));
    layer2_outputs(5113) <= not((layer1_outputs(10238)) or (layer1_outputs(8827)));
    layer2_outputs(5114) <= not(layer1_outputs(7948));
    layer2_outputs(5115) <= layer1_outputs(7162);
    layer2_outputs(5116) <= not(layer1_outputs(2126));
    layer2_outputs(5117) <= not(layer1_outputs(4588)) or (layer1_outputs(6578));
    layer2_outputs(5118) <= not(layer1_outputs(2843));
    layer2_outputs(5119) <= not(layer1_outputs(2938));
    layer2_outputs(5120) <= not(layer1_outputs(7893));
    layer2_outputs(5121) <= not(layer1_outputs(3293));
    layer2_outputs(5122) <= layer1_outputs(2325);
    layer2_outputs(5123) <= (layer1_outputs(4129)) or (layer1_outputs(6199));
    layer2_outputs(5124) <= not((layer1_outputs(5336)) xor (layer1_outputs(6685)));
    layer2_outputs(5125) <= (layer1_outputs(4333)) xor (layer1_outputs(3359));
    layer2_outputs(5126) <= not((layer1_outputs(9864)) and (layer1_outputs(468)));
    layer2_outputs(5127) <= (layer1_outputs(4594)) and (layer1_outputs(1663));
    layer2_outputs(5128) <= not((layer1_outputs(5521)) or (layer1_outputs(4533)));
    layer2_outputs(5129) <= not(layer1_outputs(937));
    layer2_outputs(5130) <= (layer1_outputs(6673)) or (layer1_outputs(1590));
    layer2_outputs(5131) <= (layer1_outputs(598)) or (layer1_outputs(2146));
    layer2_outputs(5132) <= (layer1_outputs(9400)) xor (layer1_outputs(3367));
    layer2_outputs(5133) <= (layer1_outputs(3546)) and not (layer1_outputs(2047));
    layer2_outputs(5134) <= layer1_outputs(5164);
    layer2_outputs(5135) <= not(layer1_outputs(85));
    layer2_outputs(5136) <= not(layer1_outputs(9531));
    layer2_outputs(5137) <= (layer1_outputs(2533)) xor (layer1_outputs(1445));
    layer2_outputs(5138) <= not(layer1_outputs(1575));
    layer2_outputs(5139) <= not(layer1_outputs(4791));
    layer2_outputs(5140) <= not(layer1_outputs(2100)) or (layer1_outputs(9386));
    layer2_outputs(5141) <= not(layer1_outputs(7788));
    layer2_outputs(5142) <= layer1_outputs(8660);
    layer2_outputs(5143) <= (layer1_outputs(5984)) xor (layer1_outputs(8299));
    layer2_outputs(5144) <= (layer1_outputs(1145)) and not (layer1_outputs(7402));
    layer2_outputs(5145) <= not((layer1_outputs(10010)) or (layer1_outputs(5128)));
    layer2_outputs(5146) <= (layer1_outputs(7804)) and (layer1_outputs(7729));
    layer2_outputs(5147) <= not((layer1_outputs(8842)) or (layer1_outputs(9186)));
    layer2_outputs(5148) <= layer1_outputs(7817);
    layer2_outputs(5149) <= layer1_outputs(6452);
    layer2_outputs(5150) <= not(layer1_outputs(7449)) or (layer1_outputs(5492));
    layer2_outputs(5151) <= layer1_outputs(3544);
    layer2_outputs(5152) <= layer1_outputs(5284);
    layer2_outputs(5153) <= not((layer1_outputs(4434)) and (layer1_outputs(5260)));
    layer2_outputs(5154) <= (layer1_outputs(9109)) xor (layer1_outputs(8519));
    layer2_outputs(5155) <= not(layer1_outputs(237));
    layer2_outputs(5156) <= not((layer1_outputs(4738)) and (layer1_outputs(5871)));
    layer2_outputs(5157) <= not(layer1_outputs(5087)) or (layer1_outputs(4814));
    layer2_outputs(5158) <= not((layer1_outputs(7722)) or (layer1_outputs(2597)));
    layer2_outputs(5159) <= not(layer1_outputs(7306)) or (layer1_outputs(9055));
    layer2_outputs(5160) <= not((layer1_outputs(4819)) or (layer1_outputs(5887)));
    layer2_outputs(5161) <= not(layer1_outputs(5744)) or (layer1_outputs(9778));
    layer2_outputs(5162) <= not((layer1_outputs(2147)) and (layer1_outputs(9547)));
    layer2_outputs(5163) <= layer1_outputs(7327);
    layer2_outputs(5164) <= layer1_outputs(9386);
    layer2_outputs(5165) <= (layer1_outputs(4026)) and not (layer1_outputs(7093));
    layer2_outputs(5166) <= layer1_outputs(8732);
    layer2_outputs(5167) <= not(layer1_outputs(6694));
    layer2_outputs(5168) <= (layer1_outputs(8082)) and (layer1_outputs(4080));
    layer2_outputs(5169) <= layer1_outputs(4526);
    layer2_outputs(5170) <= layer1_outputs(9586);
    layer2_outputs(5171) <= (layer1_outputs(1782)) and not (layer1_outputs(4150));
    layer2_outputs(5172) <= not(layer1_outputs(2987)) or (layer1_outputs(4567));
    layer2_outputs(5173) <= not(layer1_outputs(5921));
    layer2_outputs(5174) <= layer1_outputs(7079);
    layer2_outputs(5175) <= not(layer1_outputs(213));
    layer2_outputs(5176) <= not(layer1_outputs(1046)) or (layer1_outputs(904));
    layer2_outputs(5177) <= not((layer1_outputs(3327)) xor (layer1_outputs(3992)));
    layer2_outputs(5178) <= not(layer1_outputs(5257));
    layer2_outputs(5179) <= not((layer1_outputs(5072)) and (layer1_outputs(2788)));
    layer2_outputs(5180) <= layer1_outputs(6067);
    layer2_outputs(5181) <= not(layer1_outputs(2668));
    layer2_outputs(5182) <= not((layer1_outputs(5101)) or (layer1_outputs(7942)));
    layer2_outputs(5183) <= (layer1_outputs(9932)) xor (layer1_outputs(7438));
    layer2_outputs(5184) <= (layer1_outputs(3045)) and not (layer1_outputs(1790));
    layer2_outputs(5185) <= not(layer1_outputs(7732));
    layer2_outputs(5186) <= (layer1_outputs(6172)) or (layer1_outputs(5850));
    layer2_outputs(5187) <= (layer1_outputs(7920)) and not (layer1_outputs(2950));
    layer2_outputs(5188) <= layer1_outputs(7029);
    layer2_outputs(5189) <= layer1_outputs(6069);
    layer2_outputs(5190) <= '1';
    layer2_outputs(5191) <= (layer1_outputs(2810)) or (layer1_outputs(3031));
    layer2_outputs(5192) <= (layer1_outputs(2276)) or (layer1_outputs(9983));
    layer2_outputs(5193) <= not(layer1_outputs(8909)) or (layer1_outputs(4585));
    layer2_outputs(5194) <= (layer1_outputs(5497)) and (layer1_outputs(7234));
    layer2_outputs(5195) <= not((layer1_outputs(5064)) and (layer1_outputs(7627)));
    layer2_outputs(5196) <= (layer1_outputs(8832)) and not (layer1_outputs(7746));
    layer2_outputs(5197) <= not(layer1_outputs(3011)) or (layer1_outputs(2288));
    layer2_outputs(5198) <= not(layer1_outputs(4631));
    layer2_outputs(5199) <= not(layer1_outputs(999));
    layer2_outputs(5200) <= not(layer1_outputs(1478));
    layer2_outputs(5201) <= (layer1_outputs(4316)) and (layer1_outputs(987));
    layer2_outputs(5202) <= '1';
    layer2_outputs(5203) <= not(layer1_outputs(2879));
    layer2_outputs(5204) <= (layer1_outputs(4555)) and not (layer1_outputs(4843));
    layer2_outputs(5205) <= layer1_outputs(6941);
    layer2_outputs(5206) <= not((layer1_outputs(8350)) and (layer1_outputs(3744)));
    layer2_outputs(5207) <= not((layer1_outputs(4015)) xor (layer1_outputs(8309)));
    layer2_outputs(5208) <= layer1_outputs(8502);
    layer2_outputs(5209) <= not(layer1_outputs(3092));
    layer2_outputs(5210) <= (layer1_outputs(7553)) or (layer1_outputs(8122));
    layer2_outputs(5211) <= (layer1_outputs(6973)) and not (layer1_outputs(6250));
    layer2_outputs(5212) <= not(layer1_outputs(5622)) or (layer1_outputs(3076));
    layer2_outputs(5213) <= layer1_outputs(857);
    layer2_outputs(5214) <= not(layer1_outputs(8472)) or (layer1_outputs(7396));
    layer2_outputs(5215) <= not(layer1_outputs(9954));
    layer2_outputs(5216) <= layer1_outputs(7601);
    layer2_outputs(5217) <= not(layer1_outputs(1905));
    layer2_outputs(5218) <= not(layer1_outputs(5192)) or (layer1_outputs(1358));
    layer2_outputs(5219) <= (layer1_outputs(5516)) and not (layer1_outputs(287));
    layer2_outputs(5220) <= not((layer1_outputs(5217)) or (layer1_outputs(9020)));
    layer2_outputs(5221) <= (layer1_outputs(225)) and not (layer1_outputs(1565));
    layer2_outputs(5222) <= not(layer1_outputs(4926)) or (layer1_outputs(9117));
    layer2_outputs(5223) <= layer1_outputs(1355);
    layer2_outputs(5224) <= not(layer1_outputs(2198));
    layer2_outputs(5225) <= not((layer1_outputs(3588)) or (layer1_outputs(6197)));
    layer2_outputs(5226) <= not((layer1_outputs(7936)) xor (layer1_outputs(6982)));
    layer2_outputs(5227) <= layer1_outputs(10124);
    layer2_outputs(5228) <= layer1_outputs(4951);
    layer2_outputs(5229) <= layer1_outputs(5458);
    layer2_outputs(5230) <= (layer1_outputs(5082)) and not (layer1_outputs(7007));
    layer2_outputs(5231) <= (layer1_outputs(2456)) or (layer1_outputs(5691));
    layer2_outputs(5232) <= (layer1_outputs(1057)) or (layer1_outputs(4612));
    layer2_outputs(5233) <= not((layer1_outputs(5292)) xor (layer1_outputs(9347)));
    layer2_outputs(5234) <= (layer1_outputs(7030)) and not (layer1_outputs(1108));
    layer2_outputs(5235) <= layer1_outputs(7548);
    layer2_outputs(5236) <= not(layer1_outputs(3685));
    layer2_outputs(5237) <= not(layer1_outputs(5728)) or (layer1_outputs(7944));
    layer2_outputs(5238) <= not(layer1_outputs(8763));
    layer2_outputs(5239) <= not(layer1_outputs(9827));
    layer2_outputs(5240) <= not(layer1_outputs(3209)) or (layer1_outputs(10126));
    layer2_outputs(5241) <= layer1_outputs(296);
    layer2_outputs(5242) <= '1';
    layer2_outputs(5243) <= not(layer1_outputs(9921)) or (layer1_outputs(7368));
    layer2_outputs(5244) <= not(layer1_outputs(8924));
    layer2_outputs(5245) <= layer1_outputs(619);
    layer2_outputs(5246) <= (layer1_outputs(7482)) and (layer1_outputs(4078));
    layer2_outputs(5247) <= layer1_outputs(5360);
    layer2_outputs(5248) <= not((layer1_outputs(7437)) and (layer1_outputs(927)));
    layer2_outputs(5249) <= layer1_outputs(910);
    layer2_outputs(5250) <= (layer1_outputs(9178)) xor (layer1_outputs(8028));
    layer2_outputs(5251) <= not(layer1_outputs(5153)) or (layer1_outputs(8274));
    layer2_outputs(5252) <= not(layer1_outputs(6115));
    layer2_outputs(5253) <= not(layer1_outputs(5242));
    layer2_outputs(5254) <= (layer1_outputs(135)) xor (layer1_outputs(10147));
    layer2_outputs(5255) <= (layer1_outputs(4980)) and (layer1_outputs(3921));
    layer2_outputs(5256) <= (layer1_outputs(4210)) and not (layer1_outputs(826));
    layer2_outputs(5257) <= layer1_outputs(7319);
    layer2_outputs(5258) <= layer1_outputs(8174);
    layer2_outputs(5259) <= not(layer1_outputs(2006));
    layer2_outputs(5260) <= (layer1_outputs(7908)) or (layer1_outputs(9421));
    layer2_outputs(5261) <= not(layer1_outputs(2347));
    layer2_outputs(5262) <= not(layer1_outputs(4996)) or (layer1_outputs(2964));
    layer2_outputs(5263) <= not(layer1_outputs(9410));
    layer2_outputs(5264) <= not(layer1_outputs(968));
    layer2_outputs(5265) <= not(layer1_outputs(8292));
    layer2_outputs(5266) <= layer1_outputs(9598);
    layer2_outputs(5267) <= layer1_outputs(1554);
    layer2_outputs(5268) <= layer1_outputs(7792);
    layer2_outputs(5269) <= (layer1_outputs(4740)) xor (layer1_outputs(962));
    layer2_outputs(5270) <= (layer1_outputs(6422)) and (layer1_outputs(771));
    layer2_outputs(5271) <= not(layer1_outputs(3653));
    layer2_outputs(5272) <= (layer1_outputs(9646)) xor (layer1_outputs(8175));
    layer2_outputs(5273) <= not((layer1_outputs(4346)) xor (layer1_outputs(1103)));
    layer2_outputs(5274) <= not(layer1_outputs(8720)) or (layer1_outputs(1690));
    layer2_outputs(5275) <= not(layer1_outputs(5511));
    layer2_outputs(5276) <= layer1_outputs(9532);
    layer2_outputs(5277) <= not((layer1_outputs(5628)) and (layer1_outputs(2824)));
    layer2_outputs(5278) <= layer1_outputs(1588);
    layer2_outputs(5279) <= not(layer1_outputs(6145)) or (layer1_outputs(8068));
    layer2_outputs(5280) <= layer1_outputs(6278);
    layer2_outputs(5281) <= not(layer1_outputs(2752)) or (layer1_outputs(2798));
    layer2_outputs(5282) <= not(layer1_outputs(10209));
    layer2_outputs(5283) <= layer1_outputs(7910);
    layer2_outputs(5284) <= (layer1_outputs(6387)) xor (layer1_outputs(8330));
    layer2_outputs(5285) <= not(layer1_outputs(4659));
    layer2_outputs(5286) <= (layer1_outputs(8283)) and not (layer1_outputs(2740));
    layer2_outputs(5287) <= not((layer1_outputs(5278)) xor (layer1_outputs(8649)));
    layer2_outputs(5288) <= (layer1_outputs(9041)) xor (layer1_outputs(8861));
    layer2_outputs(5289) <= not((layer1_outputs(6130)) or (layer1_outputs(2795)));
    layer2_outputs(5290) <= not(layer1_outputs(8746));
    layer2_outputs(5291) <= not(layer1_outputs(178));
    layer2_outputs(5292) <= not((layer1_outputs(1102)) or (layer1_outputs(345)));
    layer2_outputs(5293) <= not(layer1_outputs(7322));
    layer2_outputs(5294) <= not((layer1_outputs(5245)) and (layer1_outputs(783)));
    layer2_outputs(5295) <= not(layer1_outputs(9601));
    layer2_outputs(5296) <= not((layer1_outputs(4463)) and (layer1_outputs(6852)));
    layer2_outputs(5297) <= (layer1_outputs(1199)) xor (layer1_outputs(9111));
    layer2_outputs(5298) <= (layer1_outputs(7326)) and not (layer1_outputs(4594));
    layer2_outputs(5299) <= (layer1_outputs(6236)) and not (layer1_outputs(2905));
    layer2_outputs(5300) <= not((layer1_outputs(2414)) xor (layer1_outputs(4639)));
    layer2_outputs(5301) <= not(layer1_outputs(8396));
    layer2_outputs(5302) <= (layer1_outputs(2688)) or (layer1_outputs(9149));
    layer2_outputs(5303) <= not((layer1_outputs(10071)) or (layer1_outputs(8761)));
    layer2_outputs(5304) <= not((layer1_outputs(935)) and (layer1_outputs(1326)));
    layer2_outputs(5305) <= not(layer1_outputs(6356));
    layer2_outputs(5306) <= not((layer1_outputs(6813)) and (layer1_outputs(1206)));
    layer2_outputs(5307) <= layer1_outputs(277);
    layer2_outputs(5308) <= layer1_outputs(7398);
    layer2_outputs(5309) <= (layer1_outputs(2263)) and not (layer1_outputs(142));
    layer2_outputs(5310) <= not(layer1_outputs(9453));
    layer2_outputs(5311) <= not((layer1_outputs(9755)) xor (layer1_outputs(7570)));
    layer2_outputs(5312) <= layer1_outputs(8276);
    layer2_outputs(5313) <= not(layer1_outputs(7848));
    layer2_outputs(5314) <= not(layer1_outputs(6428)) or (layer1_outputs(3547));
    layer2_outputs(5315) <= not((layer1_outputs(51)) or (layer1_outputs(4916)));
    layer2_outputs(5316) <= (layer1_outputs(9971)) and not (layer1_outputs(5373));
    layer2_outputs(5317) <= '0';
    layer2_outputs(5318) <= (layer1_outputs(6723)) and not (layer1_outputs(5337));
    layer2_outputs(5319) <= not((layer1_outputs(9179)) xor (layer1_outputs(8638)));
    layer2_outputs(5320) <= layer1_outputs(7597);
    layer2_outputs(5321) <= not(layer1_outputs(368)) or (layer1_outputs(9541));
    layer2_outputs(5322) <= not(layer1_outputs(7213));
    layer2_outputs(5323) <= layer1_outputs(8106);
    layer2_outputs(5324) <= not(layer1_outputs(1456));
    layer2_outputs(5325) <= layer1_outputs(6496);
    layer2_outputs(5326) <= not(layer1_outputs(8720));
    layer2_outputs(5327) <= not(layer1_outputs(7366));
    layer2_outputs(5328) <= not(layer1_outputs(6063));
    layer2_outputs(5329) <= not(layer1_outputs(2989)) or (layer1_outputs(902));
    layer2_outputs(5330) <= (layer1_outputs(5021)) and (layer1_outputs(9040));
    layer2_outputs(5331) <= (layer1_outputs(8322)) or (layer1_outputs(2171));
    layer2_outputs(5332) <= layer1_outputs(2419);
    layer2_outputs(5333) <= not(layer1_outputs(3543)) or (layer1_outputs(2999));
    layer2_outputs(5334) <= not(layer1_outputs(5313));
    layer2_outputs(5335) <= not((layer1_outputs(3248)) xor (layer1_outputs(8887)));
    layer2_outputs(5336) <= not(layer1_outputs(2911));
    layer2_outputs(5337) <= not(layer1_outputs(7808));
    layer2_outputs(5338) <= not(layer1_outputs(6394)) or (layer1_outputs(46));
    layer2_outputs(5339) <= not((layer1_outputs(8723)) and (layer1_outputs(8042)));
    layer2_outputs(5340) <= not((layer1_outputs(8731)) xor (layer1_outputs(7405)));
    layer2_outputs(5341) <= (layer1_outputs(6783)) xor (layer1_outputs(5103));
    layer2_outputs(5342) <= (layer1_outputs(1486)) and not (layer1_outputs(629));
    layer2_outputs(5343) <= not(layer1_outputs(9864));
    layer2_outputs(5344) <= (layer1_outputs(4021)) and (layer1_outputs(9482));
    layer2_outputs(5345) <= not(layer1_outputs(3241)) or (layer1_outputs(5394));
    layer2_outputs(5346) <= not(layer1_outputs(7058));
    layer2_outputs(5347) <= not(layer1_outputs(777)) or (layer1_outputs(7879));
    layer2_outputs(5348) <= not((layer1_outputs(2588)) and (layer1_outputs(779)));
    layer2_outputs(5349) <= not(layer1_outputs(8662)) or (layer1_outputs(7381));
    layer2_outputs(5350) <= layer1_outputs(8206);
    layer2_outputs(5351) <= layer1_outputs(6551);
    layer2_outputs(5352) <= layer1_outputs(2359);
    layer2_outputs(5353) <= layer1_outputs(140);
    layer2_outputs(5354) <= not(layer1_outputs(9602));
    layer2_outputs(5355) <= not(layer1_outputs(8569));
    layer2_outputs(5356) <= not((layer1_outputs(7584)) xor (layer1_outputs(2994)));
    layer2_outputs(5357) <= layer1_outputs(5745);
    layer2_outputs(5358) <= not(layer1_outputs(8683));
    layer2_outputs(5359) <= not(layer1_outputs(2769));
    layer2_outputs(5360) <= layer1_outputs(5982);
    layer2_outputs(5361) <= (layer1_outputs(7496)) and not (layer1_outputs(4396));
    layer2_outputs(5362) <= layer1_outputs(485);
    layer2_outputs(5363) <= (layer1_outputs(6749)) xor (layer1_outputs(7182));
    layer2_outputs(5364) <= (layer1_outputs(1812)) or (layer1_outputs(5376));
    layer2_outputs(5365) <= not((layer1_outputs(5589)) and (layer1_outputs(1543)));
    layer2_outputs(5366) <= not(layer1_outputs(9038));
    layer2_outputs(5367) <= layer1_outputs(9907);
    layer2_outputs(5368) <= (layer1_outputs(2184)) and (layer1_outputs(9605));
    layer2_outputs(5369) <= not((layer1_outputs(6435)) and (layer1_outputs(1414)));
    layer2_outputs(5370) <= (layer1_outputs(6707)) and not (layer1_outputs(5226));
    layer2_outputs(5371) <= layer1_outputs(7412);
    layer2_outputs(5372) <= (layer1_outputs(10117)) and (layer1_outputs(1351));
    layer2_outputs(5373) <= not((layer1_outputs(343)) or (layer1_outputs(2811)));
    layer2_outputs(5374) <= (layer1_outputs(7786)) or (layer1_outputs(7712));
    layer2_outputs(5375) <= layer1_outputs(9832);
    layer2_outputs(5376) <= not(layer1_outputs(1561));
    layer2_outputs(5377) <= (layer1_outputs(3497)) and not (layer1_outputs(8300));
    layer2_outputs(5378) <= not(layer1_outputs(4059)) or (layer1_outputs(8808));
    layer2_outputs(5379) <= not(layer1_outputs(5338));
    layer2_outputs(5380) <= (layer1_outputs(3364)) and not (layer1_outputs(8156));
    layer2_outputs(5381) <= (layer1_outputs(2919)) or (layer1_outputs(7333));
    layer2_outputs(5382) <= layer1_outputs(284);
    layer2_outputs(5383) <= not((layer1_outputs(10134)) xor (layer1_outputs(5544)));
    layer2_outputs(5384) <= not(layer1_outputs(6426));
    layer2_outputs(5385) <= (layer1_outputs(6227)) and (layer1_outputs(3783));
    layer2_outputs(5386) <= (layer1_outputs(1754)) and (layer1_outputs(8322));
    layer2_outputs(5387) <= not((layer1_outputs(2756)) xor (layer1_outputs(5100)));
    layer2_outputs(5388) <= layer1_outputs(6787);
    layer2_outputs(5389) <= not((layer1_outputs(9232)) and (layer1_outputs(7254)));
    layer2_outputs(5390) <= not(layer1_outputs(4050));
    layer2_outputs(5391) <= not(layer1_outputs(5839));
    layer2_outputs(5392) <= not(layer1_outputs(6329));
    layer2_outputs(5393) <= (layer1_outputs(10112)) and not (layer1_outputs(5206));
    layer2_outputs(5394) <= not((layer1_outputs(3535)) or (layer1_outputs(4074)));
    layer2_outputs(5395) <= (layer1_outputs(7399)) xor (layer1_outputs(3772));
    layer2_outputs(5396) <= (layer1_outputs(1226)) and not (layer1_outputs(2459));
    layer2_outputs(5397) <= not(layer1_outputs(5729));
    layer2_outputs(5398) <= not((layer1_outputs(6975)) xor (layer1_outputs(7874)));
    layer2_outputs(5399) <= layer1_outputs(2081);
    layer2_outputs(5400) <= not((layer1_outputs(1247)) and (layer1_outputs(9456)));
    layer2_outputs(5401) <= not(layer1_outputs(5460)) or (layer1_outputs(7041));
    layer2_outputs(5402) <= (layer1_outputs(8399)) and not (layer1_outputs(6042));
    layer2_outputs(5403) <= not(layer1_outputs(4916));
    layer2_outputs(5404) <= not(layer1_outputs(5636));
    layer2_outputs(5405) <= (layer1_outputs(8415)) or (layer1_outputs(8874));
    layer2_outputs(5406) <= not((layer1_outputs(8903)) or (layer1_outputs(6096)));
    layer2_outputs(5407) <= (layer1_outputs(6041)) xor (layer1_outputs(141));
    layer2_outputs(5408) <= not((layer1_outputs(202)) or (layer1_outputs(3393)));
    layer2_outputs(5409) <= layer1_outputs(3655);
    layer2_outputs(5410) <= (layer1_outputs(3441)) xor (layer1_outputs(1287));
    layer2_outputs(5411) <= not(layer1_outputs(6776));
    layer2_outputs(5412) <= layer1_outputs(5723);
    layer2_outputs(5413) <= not(layer1_outputs(5684)) or (layer1_outputs(8082));
    layer2_outputs(5414) <= not((layer1_outputs(7417)) or (layer1_outputs(2431)));
    layer2_outputs(5415) <= layer1_outputs(10059);
    layer2_outputs(5416) <= layer1_outputs(7736);
    layer2_outputs(5417) <= layer1_outputs(7433);
    layer2_outputs(5418) <= not(layer1_outputs(2630));
    layer2_outputs(5419) <= not(layer1_outputs(3373)) or (layer1_outputs(7947));
    layer2_outputs(5420) <= not(layer1_outputs(5695));
    layer2_outputs(5421) <= (layer1_outputs(8107)) and (layer1_outputs(5630));
    layer2_outputs(5422) <= not(layer1_outputs(33));
    layer2_outputs(5423) <= not(layer1_outputs(3658));
    layer2_outputs(5424) <= not((layer1_outputs(5765)) and (layer1_outputs(6657)));
    layer2_outputs(5425) <= not((layer1_outputs(8025)) or (layer1_outputs(4708)));
    layer2_outputs(5426) <= not(layer1_outputs(8384));
    layer2_outputs(5427) <= '1';
    layer2_outputs(5428) <= not(layer1_outputs(1007));
    layer2_outputs(5429) <= not(layer1_outputs(4125));
    layer2_outputs(5430) <= layer1_outputs(7115);
    layer2_outputs(5431) <= layer1_outputs(8857);
    layer2_outputs(5432) <= (layer1_outputs(2749)) and not (layer1_outputs(3540));
    layer2_outputs(5433) <= layer1_outputs(5496);
    layer2_outputs(5434) <= (layer1_outputs(5957)) and not (layer1_outputs(2324));
    layer2_outputs(5435) <= not(layer1_outputs(4419));
    layer2_outputs(5436) <= (layer1_outputs(5522)) and not (layer1_outputs(10050));
    layer2_outputs(5437) <= '0';
    layer2_outputs(5438) <= (layer1_outputs(6633)) and (layer1_outputs(3043));
    layer2_outputs(5439) <= (layer1_outputs(4242)) and (layer1_outputs(9074));
    layer2_outputs(5440) <= layer1_outputs(484);
    layer2_outputs(5441) <= (layer1_outputs(5775)) xor (layer1_outputs(7189));
    layer2_outputs(5442) <= not(layer1_outputs(8661)) or (layer1_outputs(1072));
    layer2_outputs(5443) <= (layer1_outputs(4367)) or (layer1_outputs(8787));
    layer2_outputs(5444) <= not(layer1_outputs(3356));
    layer2_outputs(5445) <= layer1_outputs(3115);
    layer2_outputs(5446) <= not((layer1_outputs(7035)) or (layer1_outputs(5934)));
    layer2_outputs(5447) <= (layer1_outputs(2924)) or (layer1_outputs(8842));
    layer2_outputs(5448) <= not(layer1_outputs(5615)) or (layer1_outputs(7546));
    layer2_outputs(5449) <= (layer1_outputs(3744)) and not (layer1_outputs(817));
    layer2_outputs(5450) <= (layer1_outputs(4139)) or (layer1_outputs(2363));
    layer2_outputs(5451) <= layer1_outputs(9086);
    layer2_outputs(5452) <= not(layer1_outputs(4811));
    layer2_outputs(5453) <= not(layer1_outputs(7831));
    layer2_outputs(5454) <= not(layer1_outputs(8927));
    layer2_outputs(5455) <= (layer1_outputs(4928)) and not (layer1_outputs(3992));
    layer2_outputs(5456) <= (layer1_outputs(9764)) xor (layer1_outputs(7662));
    layer2_outputs(5457) <= (layer1_outputs(1254)) or (layer1_outputs(8538));
    layer2_outputs(5458) <= not(layer1_outputs(3527));
    layer2_outputs(5459) <= (layer1_outputs(3019)) xor (layer1_outputs(4952));
    layer2_outputs(5460) <= not(layer1_outputs(5580));
    layer2_outputs(5461) <= not(layer1_outputs(5660)) or (layer1_outputs(3964));
    layer2_outputs(5462) <= not(layer1_outputs(3382));
    layer2_outputs(5463) <= (layer1_outputs(6868)) and (layer1_outputs(1613));
    layer2_outputs(5464) <= not(layer1_outputs(185));
    layer2_outputs(5465) <= not(layer1_outputs(8947));
    layer2_outputs(5466) <= not(layer1_outputs(4137)) or (layer1_outputs(1463));
    layer2_outputs(5467) <= not(layer1_outputs(9892));
    layer2_outputs(5468) <= not(layer1_outputs(5434));
    layer2_outputs(5469) <= not(layer1_outputs(9030));
    layer2_outputs(5470) <= layer1_outputs(7300);
    layer2_outputs(5471) <= layer1_outputs(2112);
    layer2_outputs(5472) <= layer1_outputs(1723);
    layer2_outputs(5473) <= (layer1_outputs(8015)) and not (layer1_outputs(639));
    layer2_outputs(5474) <= not(layer1_outputs(5151)) or (layer1_outputs(10225));
    layer2_outputs(5475) <= (layer1_outputs(2974)) and not (layer1_outputs(648));
    layer2_outputs(5476) <= layer1_outputs(6595);
    layer2_outputs(5477) <= not((layer1_outputs(3866)) or (layer1_outputs(3453)));
    layer2_outputs(5478) <= not(layer1_outputs(4247));
    layer2_outputs(5479) <= (layer1_outputs(980)) xor (layer1_outputs(7170));
    layer2_outputs(5480) <= layer1_outputs(8845);
    layer2_outputs(5481) <= not(layer1_outputs(8684));
    layer2_outputs(5482) <= not(layer1_outputs(1428));
    layer2_outputs(5483) <= layer1_outputs(4829);
    layer2_outputs(5484) <= not((layer1_outputs(803)) xor (layer1_outputs(8544)));
    layer2_outputs(5485) <= not((layer1_outputs(7121)) or (layer1_outputs(6389)));
    layer2_outputs(5486) <= layer1_outputs(5814);
    layer2_outputs(5487) <= layer1_outputs(10193);
    layer2_outputs(5488) <= not(layer1_outputs(9500)) or (layer1_outputs(3869));
    layer2_outputs(5489) <= not(layer1_outputs(304)) or (layer1_outputs(5405));
    layer2_outputs(5490) <= (layer1_outputs(1081)) and not (layer1_outputs(9745));
    layer2_outputs(5491) <= not(layer1_outputs(9395));
    layer2_outputs(5492) <= not(layer1_outputs(5253)) or (layer1_outputs(7054));
    layer2_outputs(5493) <= not(layer1_outputs(7699));
    layer2_outputs(5494) <= layer1_outputs(2153);
    layer2_outputs(5495) <= not(layer1_outputs(4258));
    layer2_outputs(5496) <= not(layer1_outputs(991));
    layer2_outputs(5497) <= not(layer1_outputs(3196));
    layer2_outputs(5498) <= not(layer1_outputs(9510)) or (layer1_outputs(3894));
    layer2_outputs(5499) <= not((layer1_outputs(7581)) or (layer1_outputs(6722)));
    layer2_outputs(5500) <= not(layer1_outputs(2969));
    layer2_outputs(5501) <= (layer1_outputs(6821)) xor (layer1_outputs(4108));
    layer2_outputs(5502) <= not(layer1_outputs(6350)) or (layer1_outputs(8005));
    layer2_outputs(5503) <= (layer1_outputs(4989)) and (layer1_outputs(5889));
    layer2_outputs(5504) <= layer1_outputs(7743);
    layer2_outputs(5505) <= not(layer1_outputs(6788));
    layer2_outputs(5506) <= layer1_outputs(4238);
    layer2_outputs(5507) <= layer1_outputs(5390);
    layer2_outputs(5508) <= not(layer1_outputs(1421));
    layer2_outputs(5509) <= (layer1_outputs(5266)) and (layer1_outputs(5290));
    layer2_outputs(5510) <= not(layer1_outputs(3231));
    layer2_outputs(5511) <= not(layer1_outputs(3435));
    layer2_outputs(5512) <= not(layer1_outputs(4419));
    layer2_outputs(5513) <= not(layer1_outputs(2868));
    layer2_outputs(5514) <= not((layer1_outputs(234)) xor (layer1_outputs(10008)));
    layer2_outputs(5515) <= not(layer1_outputs(1040));
    layer2_outputs(5516) <= (layer1_outputs(8164)) or (layer1_outputs(7538));
    layer2_outputs(5517) <= not(layer1_outputs(6148)) or (layer1_outputs(975));
    layer2_outputs(5518) <= not(layer1_outputs(6239));
    layer2_outputs(5519) <= layer1_outputs(3606);
    layer2_outputs(5520) <= layer1_outputs(7892);
    layer2_outputs(5521) <= (layer1_outputs(4465)) or (layer1_outputs(2847));
    layer2_outputs(5522) <= not((layer1_outputs(5659)) or (layer1_outputs(1155)));
    layer2_outputs(5523) <= (layer1_outputs(9219)) and not (layer1_outputs(9993));
    layer2_outputs(5524) <= not((layer1_outputs(6298)) xor (layer1_outputs(6901)));
    layer2_outputs(5525) <= (layer1_outputs(7132)) and not (layer1_outputs(4770));
    layer2_outputs(5526) <= (layer1_outputs(6606)) and not (layer1_outputs(6774));
    layer2_outputs(5527) <= not(layer1_outputs(1714)) or (layer1_outputs(6187));
    layer2_outputs(5528) <= not(layer1_outputs(2286)) or (layer1_outputs(8496));
    layer2_outputs(5529) <= not(layer1_outputs(9610)) or (layer1_outputs(4707));
    layer2_outputs(5530) <= not(layer1_outputs(7223));
    layer2_outputs(5531) <= (layer1_outputs(8956)) xor (layer1_outputs(7579));
    layer2_outputs(5532) <= not(layer1_outputs(2966));
    layer2_outputs(5533) <= layer1_outputs(1528);
    layer2_outputs(5534) <= not(layer1_outputs(1374));
    layer2_outputs(5535) <= not(layer1_outputs(3997)) or (layer1_outputs(5625));
    layer2_outputs(5536) <= layer1_outputs(5382);
    layer2_outputs(5537) <= not((layer1_outputs(2127)) xor (layer1_outputs(6542)));
    layer2_outputs(5538) <= layer1_outputs(188);
    layer2_outputs(5539) <= (layer1_outputs(8106)) and not (layer1_outputs(8775));
    layer2_outputs(5540) <= '0';
    layer2_outputs(5541) <= not(layer1_outputs(2027));
    layer2_outputs(5542) <= (layer1_outputs(3920)) and not (layer1_outputs(2204));
    layer2_outputs(5543) <= (layer1_outputs(4914)) xor (layer1_outputs(4561));
    layer2_outputs(5544) <= (layer1_outputs(9126)) or (layer1_outputs(2010));
    layer2_outputs(5545) <= (layer1_outputs(10000)) and (layer1_outputs(542));
    layer2_outputs(5546) <= (layer1_outputs(8966)) xor (layer1_outputs(1086));
    layer2_outputs(5547) <= (layer1_outputs(1176)) and (layer1_outputs(8755));
    layer2_outputs(5548) <= (layer1_outputs(8312)) and not (layer1_outputs(3138));
    layer2_outputs(5549) <= not((layer1_outputs(9027)) or (layer1_outputs(9276)));
    layer2_outputs(5550) <= (layer1_outputs(4731)) or (layer1_outputs(8612));
    layer2_outputs(5551) <= not(layer1_outputs(7139)) or (layer1_outputs(1541));
    layer2_outputs(5552) <= (layer1_outputs(6162)) and not (layer1_outputs(5929));
    layer2_outputs(5553) <= not(layer1_outputs(3292));
    layer2_outputs(5554) <= layer1_outputs(7067);
    layer2_outputs(5555) <= layer1_outputs(1979);
    layer2_outputs(5556) <= not((layer1_outputs(9807)) and (layer1_outputs(4953)));
    layer2_outputs(5557) <= (layer1_outputs(3275)) or (layer1_outputs(9555));
    layer2_outputs(5558) <= not((layer1_outputs(2211)) xor (layer1_outputs(3778)));
    layer2_outputs(5559) <= (layer1_outputs(8043)) and (layer1_outputs(4095));
    layer2_outputs(5560) <= '1';
    layer2_outputs(5561) <= not((layer1_outputs(7026)) or (layer1_outputs(6384)));
    layer2_outputs(5562) <= not(layer1_outputs(7244));
    layer2_outputs(5563) <= not((layer1_outputs(3891)) and (layer1_outputs(1286)));
    layer2_outputs(5564) <= not(layer1_outputs(7628)) or (layer1_outputs(2624));
    layer2_outputs(5565) <= (layer1_outputs(1618)) xor (layer1_outputs(9190));
    layer2_outputs(5566) <= layer1_outputs(8497);
    layer2_outputs(5567) <= layer1_outputs(5823);
    layer2_outputs(5568) <= not(layer1_outputs(3490));
    layer2_outputs(5569) <= (layer1_outputs(4455)) or (layer1_outputs(8539));
    layer2_outputs(5570) <= not((layer1_outputs(1501)) xor (layer1_outputs(10179)));
    layer2_outputs(5571) <= not((layer1_outputs(5479)) xor (layer1_outputs(2903)));
    layer2_outputs(5572) <= (layer1_outputs(9414)) or (layer1_outputs(6937));
    layer2_outputs(5573) <= not(layer1_outputs(8390));
    layer2_outputs(5574) <= layer1_outputs(4258);
    layer2_outputs(5575) <= not(layer1_outputs(8268));
    layer2_outputs(5576) <= not((layer1_outputs(8429)) or (layer1_outputs(876)));
    layer2_outputs(5577) <= (layer1_outputs(4079)) or (layer1_outputs(5105));
    layer2_outputs(5578) <= layer1_outputs(2711);
    layer2_outputs(5579) <= layer1_outputs(105);
    layer2_outputs(5580) <= (layer1_outputs(9156)) xor (layer1_outputs(1022));
    layer2_outputs(5581) <= layer1_outputs(8640);
    layer2_outputs(5582) <= layer1_outputs(9702);
    layer2_outputs(5583) <= (layer1_outputs(78)) and not (layer1_outputs(6630));
    layer2_outputs(5584) <= not(layer1_outputs(4866)) or (layer1_outputs(614));
    layer2_outputs(5585) <= not(layer1_outputs(8537));
    layer2_outputs(5586) <= layer1_outputs(4659);
    layer2_outputs(5587) <= not((layer1_outputs(7811)) and (layer1_outputs(9466)));
    layer2_outputs(5588) <= (layer1_outputs(5483)) or (layer1_outputs(2718));
    layer2_outputs(5589) <= layer1_outputs(2350);
    layer2_outputs(5590) <= not(layer1_outputs(6816));
    layer2_outputs(5591) <= not(layer1_outputs(6299)) or (layer1_outputs(9880));
    layer2_outputs(5592) <= not(layer1_outputs(2936)) or (layer1_outputs(6823));
    layer2_outputs(5593) <= not(layer1_outputs(1648)) or (layer1_outputs(9461));
    layer2_outputs(5594) <= '0';
    layer2_outputs(5595) <= layer1_outputs(255);
    layer2_outputs(5596) <= not(layer1_outputs(6470));
    layer2_outputs(5597) <= layer1_outputs(5552);
    layer2_outputs(5598) <= not((layer1_outputs(5526)) or (layer1_outputs(7815)));
    layer2_outputs(5599) <= (layer1_outputs(8219)) and (layer1_outputs(4756));
    layer2_outputs(5600) <= not((layer1_outputs(7127)) or (layer1_outputs(3452)));
    layer2_outputs(5601) <= not((layer1_outputs(4278)) and (layer1_outputs(2444)));
    layer2_outputs(5602) <= not(layer1_outputs(5160));
    layer2_outputs(5603) <= not(layer1_outputs(9774)) or (layer1_outputs(1284));
    layer2_outputs(5604) <= not(layer1_outputs(8412));
    layer2_outputs(5605) <= not(layer1_outputs(9113)) or (layer1_outputs(4787));
    layer2_outputs(5606) <= not(layer1_outputs(8577)) or (layer1_outputs(8341));
    layer2_outputs(5607) <= (layer1_outputs(4236)) and not (layer1_outputs(7632));
    layer2_outputs(5608) <= (layer1_outputs(5512)) and (layer1_outputs(8375));
    layer2_outputs(5609) <= not(layer1_outputs(4058));
    layer2_outputs(5610) <= (layer1_outputs(6549)) xor (layer1_outputs(1517));
    layer2_outputs(5611) <= (layer1_outputs(5450)) and not (layer1_outputs(5868));
    layer2_outputs(5612) <= not(layer1_outputs(5161));
    layer2_outputs(5613) <= layer1_outputs(8152);
    layer2_outputs(5614) <= not(layer1_outputs(27));
    layer2_outputs(5615) <= layer1_outputs(8034);
    layer2_outputs(5616) <= not(layer1_outputs(8325));
    layer2_outputs(5617) <= not((layer1_outputs(6718)) xor (layer1_outputs(7226)));
    layer2_outputs(5618) <= (layer1_outputs(99)) xor (layer1_outputs(1493));
    layer2_outputs(5619) <= not(layer1_outputs(5379));
    layer2_outputs(5620) <= not(layer1_outputs(5906));
    layer2_outputs(5621) <= not((layer1_outputs(6617)) or (layer1_outputs(2635)));
    layer2_outputs(5622) <= not(layer1_outputs(2551));
    layer2_outputs(5623) <= not((layer1_outputs(2046)) xor (layer1_outputs(6059)));
    layer2_outputs(5624) <= (layer1_outputs(6126)) and not (layer1_outputs(4968));
    layer2_outputs(5625) <= not(layer1_outputs(9635));
    layer2_outputs(5626) <= layer1_outputs(4299);
    layer2_outputs(5627) <= not((layer1_outputs(9714)) or (layer1_outputs(6468)));
    layer2_outputs(5628) <= not(layer1_outputs(1095));
    layer2_outputs(5629) <= not(layer1_outputs(7526));
    layer2_outputs(5630) <= not(layer1_outputs(5197));
    layer2_outputs(5631) <= layer1_outputs(7707);
    layer2_outputs(5632) <= layer1_outputs(5234);
    layer2_outputs(5633) <= (layer1_outputs(10224)) xor (layer1_outputs(6903));
    layer2_outputs(5634) <= not(layer1_outputs(9817)) or (layer1_outputs(9940));
    layer2_outputs(5635) <= not(layer1_outputs(1660));
    layer2_outputs(5636) <= not(layer1_outputs(9380));
    layer2_outputs(5637) <= (layer1_outputs(6805)) and (layer1_outputs(3760));
    layer2_outputs(5638) <= not(layer1_outputs(8554));
    layer2_outputs(5639) <= not(layer1_outputs(2420));
    layer2_outputs(5640) <= not((layer1_outputs(1964)) or (layer1_outputs(3095)));
    layer2_outputs(5641) <= (layer1_outputs(3460)) and not (layer1_outputs(1946));
    layer2_outputs(5642) <= layer1_outputs(9802);
    layer2_outputs(5643) <= (layer1_outputs(7726)) and (layer1_outputs(3343));
    layer2_outputs(5644) <= (layer1_outputs(4329)) and (layer1_outputs(6670));
    layer2_outputs(5645) <= layer1_outputs(7980);
    layer2_outputs(5646) <= (layer1_outputs(9926)) and not (layer1_outputs(8746));
    layer2_outputs(5647) <= not(layer1_outputs(1344));
    layer2_outputs(5648) <= not(layer1_outputs(3493));
    layer2_outputs(5649) <= not(layer1_outputs(5393));
    layer2_outputs(5650) <= layer1_outputs(1746);
    layer2_outputs(5651) <= not(layer1_outputs(782));
    layer2_outputs(5652) <= layer1_outputs(4996);
    layer2_outputs(5653) <= not((layer1_outputs(6636)) and (layer1_outputs(8410)));
    layer2_outputs(5654) <= (layer1_outputs(1677)) or (layer1_outputs(1558));
    layer2_outputs(5655) <= (layer1_outputs(9617)) and not (layer1_outputs(7419));
    layer2_outputs(5656) <= layer1_outputs(2402);
    layer2_outputs(5657) <= not(layer1_outputs(8247)) or (layer1_outputs(5214));
    layer2_outputs(5658) <= (layer1_outputs(6928)) and not (layer1_outputs(4486));
    layer2_outputs(5659) <= (layer1_outputs(5582)) xor (layer1_outputs(4790));
    layer2_outputs(5660) <= (layer1_outputs(8155)) or (layer1_outputs(2560));
    layer2_outputs(5661) <= (layer1_outputs(6968)) and not (layer1_outputs(8723));
    layer2_outputs(5662) <= (layer1_outputs(8818)) and (layer1_outputs(627));
    layer2_outputs(5663) <= (layer1_outputs(3316)) and (layer1_outputs(7262));
    layer2_outputs(5664) <= not(layer1_outputs(3869));
    layer2_outputs(5665) <= layer1_outputs(3580);
    layer2_outputs(5666) <= not(layer1_outputs(5015)) or (layer1_outputs(3526));
    layer2_outputs(5667) <= (layer1_outputs(9415)) xor (layer1_outputs(3862));
    layer2_outputs(5668) <= layer1_outputs(9485);
    layer2_outputs(5669) <= not(layer1_outputs(1214));
    layer2_outputs(5670) <= not(layer1_outputs(8576)) or (layer1_outputs(1536));
    layer2_outputs(5671) <= not(layer1_outputs(6221));
    layer2_outputs(5672) <= not((layer1_outputs(6558)) or (layer1_outputs(4445)));
    layer2_outputs(5673) <= not(layer1_outputs(2702)) or (layer1_outputs(5599));
    layer2_outputs(5674) <= not(layer1_outputs(6878));
    layer2_outputs(5675) <= layer1_outputs(4096);
    layer2_outputs(5676) <= not(layer1_outputs(265)) or (layer1_outputs(4938));
    layer2_outputs(5677) <= not((layer1_outputs(3235)) xor (layer1_outputs(6801)));
    layer2_outputs(5678) <= layer1_outputs(8427);
    layer2_outputs(5679) <= layer1_outputs(5969);
    layer2_outputs(5680) <= not(layer1_outputs(7036));
    layer2_outputs(5681) <= not((layer1_outputs(367)) and (layer1_outputs(2732)));
    layer2_outputs(5682) <= layer1_outputs(9076);
    layer2_outputs(5683) <= not(layer1_outputs(2661));
    layer2_outputs(5684) <= (layer1_outputs(8748)) or (layer1_outputs(8630));
    layer2_outputs(5685) <= (layer1_outputs(6474)) and (layer1_outputs(8144));
    layer2_outputs(5686) <= (layer1_outputs(6382)) xor (layer1_outputs(8875));
    layer2_outputs(5687) <= layer1_outputs(5974);
    layer2_outputs(5688) <= (layer1_outputs(1517)) xor (layer1_outputs(9101));
    layer2_outputs(5689) <= not((layer1_outputs(1767)) or (layer1_outputs(7424)));
    layer2_outputs(5690) <= not((layer1_outputs(1772)) or (layer1_outputs(5455)));
    layer2_outputs(5691) <= not((layer1_outputs(3041)) and (layer1_outputs(9366)));
    layer2_outputs(5692) <= (layer1_outputs(5638)) and not (layer1_outputs(5876));
    layer2_outputs(5693) <= (layer1_outputs(9699)) or (layer1_outputs(9500));
    layer2_outputs(5694) <= not(layer1_outputs(9180));
    layer2_outputs(5695) <= not(layer1_outputs(2673));
    layer2_outputs(5696) <= not(layer1_outputs(3307));
    layer2_outputs(5697) <= (layer1_outputs(701)) and not (layer1_outputs(560));
    layer2_outputs(5698) <= not((layer1_outputs(4391)) or (layer1_outputs(5046)));
    layer2_outputs(5699) <= (layer1_outputs(2639)) xor (layer1_outputs(2187));
    layer2_outputs(5700) <= not(layer1_outputs(9218));
    layer2_outputs(5701) <= not(layer1_outputs(884));
    layer2_outputs(5702) <= not((layer1_outputs(8573)) or (layer1_outputs(6011)));
    layer2_outputs(5703) <= layer1_outputs(2952);
    layer2_outputs(5704) <= layer1_outputs(2209);
    layer2_outputs(5705) <= layer1_outputs(5519);
    layer2_outputs(5706) <= not(layer1_outputs(9991));
    layer2_outputs(5707) <= not((layer1_outputs(7558)) xor (layer1_outputs(10226)));
    layer2_outputs(5708) <= (layer1_outputs(5143)) xor (layer1_outputs(9479));
    layer2_outputs(5709) <= not((layer1_outputs(2223)) and (layer1_outputs(9229)));
    layer2_outputs(5710) <= (layer1_outputs(3101)) xor (layer1_outputs(2887));
    layer2_outputs(5711) <= not((layer1_outputs(168)) or (layer1_outputs(5111)));
    layer2_outputs(5712) <= (layer1_outputs(4424)) and not (layer1_outputs(9054));
    layer2_outputs(5713) <= (layer1_outputs(6773)) and not (layer1_outputs(8051));
    layer2_outputs(5714) <= not(layer1_outputs(2119));
    layer2_outputs(5715) <= layer1_outputs(5202);
    layer2_outputs(5716) <= not(layer1_outputs(583));
    layer2_outputs(5717) <= not((layer1_outputs(3828)) and (layer1_outputs(1752)));
    layer2_outputs(5718) <= not((layer1_outputs(4108)) or (layer1_outputs(5681)));
    layer2_outputs(5719) <= layer1_outputs(8937);
    layer2_outputs(5720) <= not((layer1_outputs(6676)) xor (layer1_outputs(6721)));
    layer2_outputs(5721) <= not(layer1_outputs(8236));
    layer2_outputs(5722) <= not(layer1_outputs(5035));
    layer2_outputs(5723) <= not((layer1_outputs(4349)) xor (layer1_outputs(9199)));
    layer2_outputs(5724) <= not(layer1_outputs(6172));
    layer2_outputs(5725) <= layer1_outputs(4625);
    layer2_outputs(5726) <= not(layer1_outputs(2182)) or (layer1_outputs(6775));
    layer2_outputs(5727) <= layer1_outputs(7241);
    layer2_outputs(5728) <= not(layer1_outputs(3313));
    layer2_outputs(5729) <= (layer1_outputs(9130)) and not (layer1_outputs(8903));
    layer2_outputs(5730) <= not((layer1_outputs(2194)) xor (layer1_outputs(6697)));
    layer2_outputs(5731) <= layer1_outputs(2332);
    layer2_outputs(5732) <= not(layer1_outputs(8858));
    layer2_outputs(5733) <= not((layer1_outputs(3959)) xor (layer1_outputs(5518)));
    layer2_outputs(5734) <= not((layer1_outputs(10192)) xor (layer1_outputs(9948)));
    layer2_outputs(5735) <= not((layer1_outputs(2856)) xor (layer1_outputs(8982)));
    layer2_outputs(5736) <= (layer1_outputs(3402)) xor (layer1_outputs(7417));
    layer2_outputs(5737) <= layer1_outputs(5256);
    layer2_outputs(5738) <= not((layer1_outputs(1933)) xor (layer1_outputs(4920)));
    layer2_outputs(5739) <= not(layer1_outputs(1225));
    layer2_outputs(5740) <= (layer1_outputs(4172)) and not (layer1_outputs(4825));
    layer2_outputs(5741) <= not(layer1_outputs(7331));
    layer2_outputs(5742) <= not(layer1_outputs(7899)) or (layer1_outputs(1627));
    layer2_outputs(5743) <= (layer1_outputs(9197)) xor (layer1_outputs(9518));
    layer2_outputs(5744) <= (layer1_outputs(3617)) and (layer1_outputs(4872));
    layer2_outputs(5745) <= (layer1_outputs(3856)) xor (layer1_outputs(5081));
    layer2_outputs(5746) <= not(layer1_outputs(4439));
    layer2_outputs(5747) <= not((layer1_outputs(1276)) or (layer1_outputs(9624)));
    layer2_outputs(5748) <= layer1_outputs(5799);
    layer2_outputs(5749) <= not(layer1_outputs(7696));
    layer2_outputs(5750) <= (layer1_outputs(8046)) or (layer1_outputs(3446));
    layer2_outputs(5751) <= layer1_outputs(9998);
    layer2_outputs(5752) <= not((layer1_outputs(5641)) xor (layer1_outputs(5269)));
    layer2_outputs(5753) <= not(layer1_outputs(3936)) or (layer1_outputs(10228));
    layer2_outputs(5754) <= (layer1_outputs(3340)) and (layer1_outputs(5892));
    layer2_outputs(5755) <= (layer1_outputs(1684)) and not (layer1_outputs(6942));
    layer2_outputs(5756) <= not(layer1_outputs(5162));
    layer2_outputs(5757) <= (layer1_outputs(2683)) and (layer1_outputs(6999));
    layer2_outputs(5758) <= (layer1_outputs(3358)) and not (layer1_outputs(6107));
    layer2_outputs(5759) <= layer1_outputs(4354);
    layer2_outputs(5760) <= not(layer1_outputs(2619)) or (layer1_outputs(7453));
    layer2_outputs(5761) <= (layer1_outputs(3133)) and not (layer1_outputs(8649));
    layer2_outputs(5762) <= not(layer1_outputs(5435));
    layer2_outputs(5763) <= not(layer1_outputs(8870)) or (layer1_outputs(4754));
    layer2_outputs(5764) <= not(layer1_outputs(2365));
    layer2_outputs(5765) <= not((layer1_outputs(7003)) and (layer1_outputs(9841)));
    layer2_outputs(5766) <= not(layer1_outputs(7129));
    layer2_outputs(5767) <= not((layer1_outputs(9691)) xor (layer1_outputs(7158)));
    layer2_outputs(5768) <= not((layer1_outputs(660)) or (layer1_outputs(8532)));
    layer2_outputs(5769) <= (layer1_outputs(2556)) and not (layer1_outputs(358));
    layer2_outputs(5770) <= layer1_outputs(9277);
    layer2_outputs(5771) <= not(layer1_outputs(9231));
    layer2_outputs(5772) <= layer1_outputs(10088);
    layer2_outputs(5773) <= (layer1_outputs(6174)) or (layer1_outputs(8142));
    layer2_outputs(5774) <= not(layer1_outputs(5850));
    layer2_outputs(5775) <= (layer1_outputs(3107)) and not (layer1_outputs(8780));
    layer2_outputs(5776) <= '0';
    layer2_outputs(5777) <= (layer1_outputs(5963)) and not (layer1_outputs(978));
    layer2_outputs(5778) <= not((layer1_outputs(4016)) or (layer1_outputs(1887)));
    layer2_outputs(5779) <= not((layer1_outputs(8698)) and (layer1_outputs(3317)));
    layer2_outputs(5780) <= layer1_outputs(244);
    layer2_outputs(5781) <= (layer1_outputs(6742)) or (layer1_outputs(1792));
    layer2_outputs(5782) <= layer1_outputs(2714);
    layer2_outputs(5783) <= (layer1_outputs(4127)) and not (layer1_outputs(9459));
    layer2_outputs(5784) <= (layer1_outputs(502)) and not (layer1_outputs(4111));
    layer2_outputs(5785) <= '0';
    layer2_outputs(5786) <= not(layer1_outputs(216));
    layer2_outputs(5787) <= (layer1_outputs(1020)) xor (layer1_outputs(5130));
    layer2_outputs(5788) <= not(layer1_outputs(2437));
    layer2_outputs(5789) <= layer1_outputs(3795);
    layer2_outputs(5790) <= (layer1_outputs(6812)) xor (layer1_outputs(3518));
    layer2_outputs(5791) <= (layer1_outputs(50)) or (layer1_outputs(5712));
    layer2_outputs(5792) <= (layer1_outputs(1012)) and not (layer1_outputs(3066));
    layer2_outputs(5793) <= (layer1_outputs(8762)) and (layer1_outputs(4311));
    layer2_outputs(5794) <= layer1_outputs(3143);
    layer2_outputs(5795) <= not(layer1_outputs(7059));
    layer2_outputs(5796) <= (layer1_outputs(117)) and (layer1_outputs(8419));
    layer2_outputs(5797) <= not((layer1_outputs(4862)) and (layer1_outputs(1202)));
    layer2_outputs(5798) <= not((layer1_outputs(2184)) and (layer1_outputs(1292)));
    layer2_outputs(5799) <= layer1_outputs(1319);
    layer2_outputs(5800) <= (layer1_outputs(9959)) or (layer1_outputs(4317));
    layer2_outputs(5801) <= (layer1_outputs(4977)) xor (layer1_outputs(7710));
    layer2_outputs(5802) <= layer1_outputs(6211);
    layer2_outputs(5803) <= not(layer1_outputs(4719));
    layer2_outputs(5804) <= not((layer1_outputs(3378)) and (layer1_outputs(3002)));
    layer2_outputs(5805) <= (layer1_outputs(2935)) or (layer1_outputs(9925));
    layer2_outputs(5806) <= layer1_outputs(8059);
    layer2_outputs(5807) <= not((layer1_outputs(2842)) xor (layer1_outputs(8016)));
    layer2_outputs(5808) <= not(layer1_outputs(8966));
    layer2_outputs(5809) <= not(layer1_outputs(10018));
    layer2_outputs(5810) <= layer1_outputs(9727);
    layer2_outputs(5811) <= not(layer1_outputs(299)) or (layer1_outputs(635));
    layer2_outputs(5812) <= not(layer1_outputs(3139)) or (layer1_outputs(8764));
    layer2_outputs(5813) <= layer1_outputs(2995);
    layer2_outputs(5814) <= not(layer1_outputs(3837)) or (layer1_outputs(5664));
    layer2_outputs(5815) <= (layer1_outputs(10105)) or (layer1_outputs(4454));
    layer2_outputs(5816) <= layer1_outputs(7365);
    layer2_outputs(5817) <= not(layer1_outputs(3854)) or (layer1_outputs(1757));
    layer2_outputs(5818) <= not(layer1_outputs(10090)) or (layer1_outputs(8423));
    layer2_outputs(5819) <= (layer1_outputs(5076)) and (layer1_outputs(6203));
    layer2_outputs(5820) <= (layer1_outputs(8303)) and not (layer1_outputs(3476));
    layer2_outputs(5821) <= not((layer1_outputs(3750)) xor (layer1_outputs(4581)));
    layer2_outputs(5822) <= not((layer1_outputs(5502)) xor (layer1_outputs(2466)));
    layer2_outputs(5823) <= (layer1_outputs(7984)) and not (layer1_outputs(5936));
    layer2_outputs(5824) <= (layer1_outputs(2068)) and (layer1_outputs(2238));
    layer2_outputs(5825) <= layer1_outputs(6480);
    layer2_outputs(5826) <= (layer1_outputs(2229)) and (layer1_outputs(7083));
    layer2_outputs(5827) <= not(layer1_outputs(6808));
    layer2_outputs(5828) <= (layer1_outputs(4175)) xor (layer1_outputs(5278));
    layer2_outputs(5829) <= (layer1_outputs(2653)) and not (layer1_outputs(9373));
    layer2_outputs(5830) <= '1';
    layer2_outputs(5831) <= layer1_outputs(851);
    layer2_outputs(5832) <= not(layer1_outputs(7003));
    layer2_outputs(5833) <= (layer1_outputs(8336)) or (layer1_outputs(5271));
    layer2_outputs(5834) <= (layer1_outputs(5001)) and not (layer1_outputs(5620));
    layer2_outputs(5835) <= not((layer1_outputs(2187)) or (layer1_outputs(6042)));
    layer2_outputs(5836) <= not(layer1_outputs(9128));
    layer2_outputs(5837) <= layer1_outputs(3080);
    layer2_outputs(5838) <= not((layer1_outputs(6260)) and (layer1_outputs(1508)));
    layer2_outputs(5839) <= (layer1_outputs(8454)) and not (layer1_outputs(7630));
    layer2_outputs(5840) <= not(layer1_outputs(4805));
    layer2_outputs(5841) <= not(layer1_outputs(1231));
    layer2_outputs(5842) <= (layer1_outputs(9200)) xor (layer1_outputs(9387));
    layer2_outputs(5843) <= not(layer1_outputs(1959));
    layer2_outputs(5844) <= layer1_outputs(2880);
    layer2_outputs(5845) <= not(layer1_outputs(5966));
    layer2_outputs(5846) <= layer1_outputs(1241);
    layer2_outputs(5847) <= layer1_outputs(1944);
    layer2_outputs(5848) <= layer1_outputs(5055);
    layer2_outputs(5849) <= layer1_outputs(8930);
    layer2_outputs(5850) <= (layer1_outputs(6958)) or (layer1_outputs(5725));
    layer2_outputs(5851) <= not(layer1_outputs(5718));
    layer2_outputs(5852) <= not(layer1_outputs(10202)) or (layer1_outputs(8875));
    layer2_outputs(5853) <= not(layer1_outputs(8493));
    layer2_outputs(5854) <= layer1_outputs(3139);
    layer2_outputs(5855) <= (layer1_outputs(6810)) or (layer1_outputs(6610));
    layer2_outputs(5856) <= layer1_outputs(814);
    layer2_outputs(5857) <= not(layer1_outputs(6264)) or (layer1_outputs(3571));
    layer2_outputs(5858) <= not(layer1_outputs(1885)) or (layer1_outputs(769));
    layer2_outputs(5859) <= not(layer1_outputs(6076));
    layer2_outputs(5860) <= (layer1_outputs(7038)) and not (layer1_outputs(5213));
    layer2_outputs(5861) <= layer1_outputs(9719);
    layer2_outputs(5862) <= layer1_outputs(7866);
    layer2_outputs(5863) <= not(layer1_outputs(9172));
    layer2_outputs(5864) <= not(layer1_outputs(8715)) or (layer1_outputs(5752));
    layer2_outputs(5865) <= layer1_outputs(1165);
    layer2_outputs(5866) <= (layer1_outputs(228)) and not (layer1_outputs(8182));
    layer2_outputs(5867) <= layer1_outputs(255);
    layer2_outputs(5868) <= (layer1_outputs(1657)) or (layer1_outputs(5530));
    layer2_outputs(5869) <= not(layer1_outputs(2034));
    layer2_outputs(5870) <= not(layer1_outputs(3023));
    layer2_outputs(5871) <= not(layer1_outputs(9217));
    layer2_outputs(5872) <= not(layer1_outputs(7393));
    layer2_outputs(5873) <= (layer1_outputs(1226)) and not (layer1_outputs(5480));
    layer2_outputs(5874) <= not(layer1_outputs(1785));
    layer2_outputs(5875) <= not((layer1_outputs(8258)) or (layer1_outputs(9990)));
    layer2_outputs(5876) <= not(layer1_outputs(3307));
    layer2_outputs(5877) <= not((layer1_outputs(4151)) and (layer1_outputs(9562)));
    layer2_outputs(5878) <= not(layer1_outputs(1549));
    layer2_outputs(5879) <= (layer1_outputs(4121)) xor (layer1_outputs(5136));
    layer2_outputs(5880) <= (layer1_outputs(10157)) or (layer1_outputs(7237));
    layer2_outputs(5881) <= not(layer1_outputs(7009));
    layer2_outputs(5882) <= not(layer1_outputs(679));
    layer2_outputs(5883) <= layer1_outputs(9384);
    layer2_outputs(5884) <= (layer1_outputs(8887)) and not (layer1_outputs(4097));
    layer2_outputs(5885) <= not(layer1_outputs(6319));
    layer2_outputs(5886) <= layer1_outputs(9671);
    layer2_outputs(5887) <= not(layer1_outputs(5623)) or (layer1_outputs(2212));
    layer2_outputs(5888) <= not(layer1_outputs(893));
    layer2_outputs(5889) <= not((layer1_outputs(4948)) and (layer1_outputs(5505)));
    layer2_outputs(5890) <= not(layer1_outputs(6898)) or (layer1_outputs(9307));
    layer2_outputs(5891) <= (layer1_outputs(3394)) xor (layer1_outputs(1738));
    layer2_outputs(5892) <= layer1_outputs(1252);
    layer2_outputs(5893) <= (layer1_outputs(9424)) and not (layer1_outputs(9614));
    layer2_outputs(5894) <= not(layer1_outputs(860));
    layer2_outputs(5895) <= (layer1_outputs(8478)) and not (layer1_outputs(8591));
    layer2_outputs(5896) <= layer1_outputs(3163);
    layer2_outputs(5897) <= '0';
    layer2_outputs(5898) <= not(layer1_outputs(7276));
    layer2_outputs(5899) <= not((layer1_outputs(6357)) and (layer1_outputs(5804)));
    layer2_outputs(5900) <= not(layer1_outputs(2970));
    layer2_outputs(5901) <= layer1_outputs(3847);
    layer2_outputs(5902) <= (layer1_outputs(8771)) or (layer1_outputs(2890));
    layer2_outputs(5903) <= not((layer1_outputs(8745)) xor (layer1_outputs(6314)));
    layer2_outputs(5904) <= not(layer1_outputs(811)) or (layer1_outputs(2537));
    layer2_outputs(5905) <= layer1_outputs(4773);
    layer2_outputs(5906) <= not((layer1_outputs(4430)) xor (layer1_outputs(9867)));
    layer2_outputs(5907) <= layer1_outputs(4069);
    layer2_outputs(5908) <= '0';
    layer2_outputs(5909) <= not(layer1_outputs(5637));
    layer2_outputs(5910) <= layer1_outputs(7281);
    layer2_outputs(5911) <= not(layer1_outputs(7173));
    layer2_outputs(5912) <= (layer1_outputs(1501)) or (layer1_outputs(653));
    layer2_outputs(5913) <= (layer1_outputs(10180)) and not (layer1_outputs(10096));
    layer2_outputs(5914) <= not(layer1_outputs(5110));
    layer2_outputs(5915) <= (layer1_outputs(4030)) and not (layer1_outputs(482));
    layer2_outputs(5916) <= layer1_outputs(1883);
    layer2_outputs(5917) <= not(layer1_outputs(984));
    layer2_outputs(5918) <= not(layer1_outputs(7603));
    layer2_outputs(5919) <= not((layer1_outputs(3251)) xor (layer1_outputs(1839)));
    layer2_outputs(5920) <= not((layer1_outputs(7156)) and (layer1_outputs(2718)));
    layer2_outputs(5921) <= not((layer1_outputs(5276)) xor (layer1_outputs(8778)));
    layer2_outputs(5922) <= (layer1_outputs(6047)) or (layer1_outputs(2704));
    layer2_outputs(5923) <= not(layer1_outputs(3838)) or (layer1_outputs(3893));
    layer2_outputs(5924) <= layer1_outputs(6179);
    layer2_outputs(5925) <= not(layer1_outputs(1932));
    layer2_outputs(5926) <= not(layer1_outputs(4318));
    layer2_outputs(5927) <= not(layer1_outputs(8798));
    layer2_outputs(5928) <= (layer1_outputs(3062)) or (layer1_outputs(8038));
    layer2_outputs(5929) <= not(layer1_outputs(8694)) or (layer1_outputs(8173));
    layer2_outputs(5930) <= (layer1_outputs(1301)) and not (layer1_outputs(75));
    layer2_outputs(5931) <= (layer1_outputs(5360)) and (layer1_outputs(625));
    layer2_outputs(5932) <= layer1_outputs(8893);
    layer2_outputs(5933) <= not((layer1_outputs(1334)) and (layer1_outputs(9988)));
    layer2_outputs(5934) <= (layer1_outputs(1670)) or (layer1_outputs(9036));
    layer2_outputs(5935) <= '0';
    layer2_outputs(5936) <= not(layer1_outputs(9093));
    layer2_outputs(5937) <= not(layer1_outputs(3427));
    layer2_outputs(5938) <= (layer1_outputs(8620)) and not (layer1_outputs(949));
    layer2_outputs(5939) <= not((layer1_outputs(6070)) xor (layer1_outputs(5154)));
    layer2_outputs(5940) <= layer1_outputs(9356);
    layer2_outputs(5941) <= '1';
    layer2_outputs(5942) <= not(layer1_outputs(6799));
    layer2_outputs(5943) <= layer1_outputs(5676);
    layer2_outputs(5944) <= not(layer1_outputs(9996));
    layer2_outputs(5945) <= (layer1_outputs(3465)) and (layer1_outputs(10062));
    layer2_outputs(5946) <= (layer1_outputs(433)) and not (layer1_outputs(4853));
    layer2_outputs(5947) <= not(layer1_outputs(8727)) or (layer1_outputs(1170));
    layer2_outputs(5948) <= not(layer1_outputs(964));
    layer2_outputs(5949) <= not(layer1_outputs(1438)) or (layer1_outputs(6267));
    layer2_outputs(5950) <= not((layer1_outputs(6890)) or (layer1_outputs(3480)));
    layer2_outputs(5951) <= (layer1_outputs(8179)) xor (layer1_outputs(7589));
    layer2_outputs(5952) <= not(layer1_outputs(1125));
    layer2_outputs(5953) <= not(layer1_outputs(6032));
    layer2_outputs(5954) <= (layer1_outputs(1619)) and not (layer1_outputs(8108));
    layer2_outputs(5955) <= not(layer1_outputs(5919));
    layer2_outputs(5956) <= not(layer1_outputs(10239));
    layer2_outputs(5957) <= not(layer1_outputs(1547));
    layer2_outputs(5958) <= layer1_outputs(3222);
    layer2_outputs(5959) <= not(layer1_outputs(2279));
    layer2_outputs(5960) <= not(layer1_outputs(5665)) or (layer1_outputs(7460));
    layer2_outputs(5961) <= not(layer1_outputs(9608));
    layer2_outputs(5962) <= not((layer1_outputs(3150)) and (layer1_outputs(3513)));
    layer2_outputs(5963) <= (layer1_outputs(742)) or (layer1_outputs(6007));
    layer2_outputs(5964) <= (layer1_outputs(4062)) or (layer1_outputs(4882));
    layer2_outputs(5965) <= layer1_outputs(3661);
    layer2_outputs(5966) <= not((layer1_outputs(1291)) xor (layer1_outputs(8331)));
    layer2_outputs(5967) <= not(layer1_outputs(1317));
    layer2_outputs(5968) <= not((layer1_outputs(8695)) and (layer1_outputs(722)));
    layer2_outputs(5969) <= not(layer1_outputs(9785)) or (layer1_outputs(10168));
    layer2_outputs(5970) <= (layer1_outputs(4623)) and (layer1_outputs(7833));
    layer2_outputs(5971) <= layer1_outputs(8070);
    layer2_outputs(5972) <= not(layer1_outputs(9330)) or (layer1_outputs(1039));
    layer2_outputs(5973) <= not(layer1_outputs(5303));
    layer2_outputs(5974) <= (layer1_outputs(9129)) and not (layer1_outputs(3774));
    layer2_outputs(5975) <= not(layer1_outputs(5558));
    layer2_outputs(5976) <= not(layer1_outputs(4501));
    layer2_outputs(5977) <= not(layer1_outputs(4799)) or (layer1_outputs(1237));
    layer2_outputs(5978) <= (layer1_outputs(5987)) xor (layer1_outputs(3195));
    layer2_outputs(5979) <= (layer1_outputs(9086)) and not (layer1_outputs(150));
    layer2_outputs(5980) <= not((layer1_outputs(10205)) or (layer1_outputs(8062)));
    layer2_outputs(5981) <= not((layer1_outputs(7457)) or (layer1_outputs(3296)));
    layer2_outputs(5982) <= not((layer1_outputs(8738)) or (layer1_outputs(9348)));
    layer2_outputs(5983) <= layer1_outputs(3759);
    layer2_outputs(5984) <= (layer1_outputs(1094)) xor (layer1_outputs(4587));
    layer2_outputs(5985) <= not((layer1_outputs(389)) xor (layer1_outputs(7332)));
    layer2_outputs(5986) <= layer1_outputs(3996);
    layer2_outputs(5987) <= (layer1_outputs(3183)) xor (layer1_outputs(6131));
    layer2_outputs(5988) <= not(layer1_outputs(7700));
    layer2_outputs(5989) <= (layer1_outputs(6236)) and (layer1_outputs(7647));
    layer2_outputs(5990) <= not(layer1_outputs(8775));
    layer2_outputs(5991) <= layer1_outputs(9971);
    layer2_outputs(5992) <= not((layer1_outputs(8895)) xor (layer1_outputs(1653)));
    layer2_outputs(5993) <= not((layer1_outputs(4147)) and (layer1_outputs(1773)));
    layer2_outputs(5994) <= (layer1_outputs(10164)) xor (layer1_outputs(3827));
    layer2_outputs(5995) <= (layer1_outputs(8944)) and not (layer1_outputs(1631));
    layer2_outputs(5996) <= not((layer1_outputs(6364)) and (layer1_outputs(4469)));
    layer2_outputs(5997) <= (layer1_outputs(8349)) and (layer1_outputs(3745));
    layer2_outputs(5998) <= (layer1_outputs(1605)) or (layer1_outputs(8057));
    layer2_outputs(5999) <= layer1_outputs(211);
    layer2_outputs(6000) <= not((layer1_outputs(5048)) and (layer1_outputs(4808)));
    layer2_outputs(6001) <= layer1_outputs(4345);
    layer2_outputs(6002) <= not((layer1_outputs(5666)) and (layer1_outputs(599)));
    layer2_outputs(6003) <= layer1_outputs(785);
    layer2_outputs(6004) <= '0';
    layer2_outputs(6005) <= layer1_outputs(7156);
    layer2_outputs(6006) <= not(layer1_outputs(695));
    layer2_outputs(6007) <= not(layer1_outputs(4863));
    layer2_outputs(6008) <= layer1_outputs(7538);
    layer2_outputs(6009) <= (layer1_outputs(9787)) and not (layer1_outputs(6284));
    layer2_outputs(6010) <= not(layer1_outputs(7470));
    layer2_outputs(6011) <= layer1_outputs(9232);
    layer2_outputs(6012) <= (layer1_outputs(3656)) or (layer1_outputs(5761));
    layer2_outputs(6013) <= not(layer1_outputs(5671));
    layer2_outputs(6014) <= layer1_outputs(9127);
    layer2_outputs(6015) <= layer1_outputs(22);
    layer2_outputs(6016) <= layer1_outputs(3653);
    layer2_outputs(6017) <= (layer1_outputs(5632)) and not (layer1_outputs(276));
    layer2_outputs(6018) <= (layer1_outputs(4206)) or (layer1_outputs(10002));
    layer2_outputs(6019) <= not((layer1_outputs(1243)) or (layer1_outputs(5082)));
    layer2_outputs(6020) <= not((layer1_outputs(8508)) xor (layer1_outputs(7962)));
    layer2_outputs(6021) <= (layer1_outputs(7184)) xor (layer1_outputs(4666));
    layer2_outputs(6022) <= layer1_outputs(5056);
    layer2_outputs(6023) <= (layer1_outputs(8990)) and not (layer1_outputs(9618));
    layer2_outputs(6024) <= (layer1_outputs(552)) or (layer1_outputs(9310));
    layer2_outputs(6025) <= (layer1_outputs(3801)) and (layer1_outputs(5446));
    layer2_outputs(6026) <= (layer1_outputs(7758)) and not (layer1_outputs(8573));
    layer2_outputs(6027) <= layer1_outputs(8593);
    layer2_outputs(6028) <= not((layer1_outputs(9263)) xor (layer1_outputs(10118)));
    layer2_outputs(6029) <= not(layer1_outputs(6780));
    layer2_outputs(6030) <= not(layer1_outputs(6153)) or (layer1_outputs(7425));
    layer2_outputs(6031) <= (layer1_outputs(601)) and not (layer1_outputs(2229));
    layer2_outputs(6032) <= (layer1_outputs(7109)) and (layer1_outputs(6866));
    layer2_outputs(6033) <= not(layer1_outputs(4937));
    layer2_outputs(6034) <= layer1_outputs(673);
    layer2_outputs(6035) <= layer1_outputs(5970);
    layer2_outputs(6036) <= layer1_outputs(7020);
    layer2_outputs(6037) <= layer1_outputs(6306);
    layer2_outputs(6038) <= not(layer1_outputs(8207));
    layer2_outputs(6039) <= not(layer1_outputs(1632)) or (layer1_outputs(8443));
    layer2_outputs(6040) <= (layer1_outputs(8920)) or (layer1_outputs(676));
    layer2_outputs(6041) <= layer1_outputs(210);
    layer2_outputs(6042) <= layer1_outputs(4241);
    layer2_outputs(6043) <= (layer1_outputs(10132)) and not (layer1_outputs(8135));
    layer2_outputs(6044) <= not(layer1_outputs(6252));
    layer2_outputs(6045) <= layer1_outputs(5754);
    layer2_outputs(6046) <= (layer1_outputs(6598)) xor (layer1_outputs(6755));
    layer2_outputs(6047) <= layer1_outputs(711);
    layer2_outputs(6048) <= layer1_outputs(10237);
    layer2_outputs(6049) <= not(layer1_outputs(6671));
    layer2_outputs(6050) <= not(layer1_outputs(4128)) or (layer1_outputs(403));
    layer2_outputs(6051) <= (layer1_outputs(5575)) and not (layer1_outputs(1096));
    layer2_outputs(6052) <= not((layer1_outputs(5002)) xor (layer1_outputs(6882)));
    layer2_outputs(6053) <= (layer1_outputs(9736)) or (layer1_outputs(9353));
    layer2_outputs(6054) <= not((layer1_outputs(8951)) and (layer1_outputs(115)));
    layer2_outputs(6055) <= (layer1_outputs(2306)) and not (layer1_outputs(209));
    layer2_outputs(6056) <= (layer1_outputs(95)) and (layer1_outputs(2075));
    layer2_outputs(6057) <= (layer1_outputs(5600)) xor (layer1_outputs(2884));
    layer2_outputs(6058) <= not(layer1_outputs(6286));
    layer2_outputs(6059) <= (layer1_outputs(5743)) and not (layer1_outputs(9678));
    layer2_outputs(6060) <= layer1_outputs(8250);
    layer2_outputs(6061) <= (layer1_outputs(6183)) and not (layer1_outputs(7936));
    layer2_outputs(6062) <= not((layer1_outputs(3823)) or (layer1_outputs(9281)));
    layer2_outputs(6063) <= not((layer1_outputs(976)) xor (layer1_outputs(2634)));
    layer2_outputs(6064) <= not((layer1_outputs(3723)) or (layer1_outputs(1256)));
    layer2_outputs(6065) <= layer1_outputs(8776);
    layer2_outputs(6066) <= not((layer1_outputs(5000)) or (layer1_outputs(5855)));
    layer2_outputs(6067) <= not(layer1_outputs(4204));
    layer2_outputs(6068) <= not(layer1_outputs(6571));
    layer2_outputs(6069) <= not(layer1_outputs(10222));
    layer2_outputs(6070) <= layer1_outputs(3602);
    layer2_outputs(6071) <= not(layer1_outputs(7462)) or (layer1_outputs(7112));
    layer2_outputs(6072) <= not(layer1_outputs(5945));
    layer2_outputs(6073) <= not(layer1_outputs(129));
    layer2_outputs(6074) <= not(layer1_outputs(6899));
    layer2_outputs(6075) <= not(layer1_outputs(9062)) or (layer1_outputs(691));
    layer2_outputs(6076) <= (layer1_outputs(8387)) xor (layer1_outputs(4634));
    layer2_outputs(6077) <= (layer1_outputs(1490)) xor (layer1_outputs(1413));
    layer2_outputs(6078) <= layer1_outputs(953);
    layer2_outputs(6079) <= not(layer1_outputs(4559));
    layer2_outputs(6080) <= (layer1_outputs(6567)) xor (layer1_outputs(7258));
    layer2_outputs(6081) <= not((layer1_outputs(8035)) or (layer1_outputs(8739)));
    layer2_outputs(6082) <= (layer1_outputs(2153)) and not (layer1_outputs(5071));
    layer2_outputs(6083) <= (layer1_outputs(5188)) or (layer1_outputs(4338));
    layer2_outputs(6084) <= (layer1_outputs(7914)) xor (layer1_outputs(9161));
    layer2_outputs(6085) <= not(layer1_outputs(6049));
    layer2_outputs(6086) <= not((layer1_outputs(3261)) xor (layer1_outputs(3728)));
    layer2_outputs(6087) <= not(layer1_outputs(29));
    layer2_outputs(6088) <= layer1_outputs(1635);
    layer2_outputs(6089) <= not((layer1_outputs(2645)) or (layer1_outputs(9676)));
    layer2_outputs(6090) <= layer1_outputs(3633);
    layer2_outputs(6091) <= (layer1_outputs(7867)) xor (layer1_outputs(2721));
    layer2_outputs(6092) <= layer1_outputs(1458);
    layer2_outputs(6093) <= not((layer1_outputs(3670)) xor (layer1_outputs(1271)));
    layer2_outputs(6094) <= not(layer1_outputs(2090)) or (layer1_outputs(751));
    layer2_outputs(6095) <= not(layer1_outputs(8568));
    layer2_outputs(6096) <= not(layer1_outputs(318));
    layer2_outputs(6097) <= (layer1_outputs(7537)) and not (layer1_outputs(8197));
    layer2_outputs(6098) <= not(layer1_outputs(7177));
    layer2_outputs(6099) <= (layer1_outputs(4214)) and (layer1_outputs(6738));
    layer2_outputs(6100) <= not((layer1_outputs(4117)) xor (layer1_outputs(1624)));
    layer2_outputs(6101) <= layer1_outputs(4900);
    layer2_outputs(6102) <= (layer1_outputs(1912)) xor (layer1_outputs(3185));
    layer2_outputs(6103) <= not(layer1_outputs(218));
    layer2_outputs(6104) <= not((layer1_outputs(5446)) xor (layer1_outputs(2447)));
    layer2_outputs(6105) <= layer1_outputs(999);
    layer2_outputs(6106) <= (layer1_outputs(1302)) xor (layer1_outputs(9396));
    layer2_outputs(6107) <= not(layer1_outputs(9878));
    layer2_outputs(6108) <= (layer1_outputs(7923)) xor (layer1_outputs(2308));
    layer2_outputs(6109) <= not(layer1_outputs(7991));
    layer2_outputs(6110) <= (layer1_outputs(5940)) and not (layer1_outputs(4915));
    layer2_outputs(6111) <= layer1_outputs(3027);
    layer2_outputs(6112) <= not((layer1_outputs(9278)) xor (layer1_outputs(9163)));
    layer2_outputs(6113) <= not(layer1_outputs(8371));
    layer2_outputs(6114) <= not(layer1_outputs(9524));
    layer2_outputs(6115) <= (layer1_outputs(3552)) and not (layer1_outputs(10102));
    layer2_outputs(6116) <= layer1_outputs(192);
    layer2_outputs(6117) <= layer1_outputs(8235);
    layer2_outputs(6118) <= not(layer1_outputs(9584));
    layer2_outputs(6119) <= layer1_outputs(6597);
    layer2_outputs(6120) <= (layer1_outputs(2839)) or (layer1_outputs(3109));
    layer2_outputs(6121) <= not(layer1_outputs(3553));
    layer2_outputs(6122) <= (layer1_outputs(8017)) and (layer1_outputs(8734));
    layer2_outputs(6123) <= layer1_outputs(2705);
    layer2_outputs(6124) <= layer1_outputs(3123);
    layer2_outputs(6125) <= layer1_outputs(3632);
    layer2_outputs(6126) <= (layer1_outputs(5028)) or (layer1_outputs(1073));
    layer2_outputs(6127) <= not((layer1_outputs(6570)) and (layer1_outputs(7990)));
    layer2_outputs(6128) <= (layer1_outputs(5841)) or (layer1_outputs(3536));
    layer2_outputs(6129) <= not(layer1_outputs(6077));
    layer2_outputs(6130) <= not(layer1_outputs(4167));
    layer2_outputs(6131) <= layer1_outputs(2608);
    layer2_outputs(6132) <= layer1_outputs(7289);
    layer2_outputs(6133) <= (layer1_outputs(5323)) or (layer1_outputs(1123));
    layer2_outputs(6134) <= (layer1_outputs(3847)) and not (layer1_outputs(4457));
    layer2_outputs(6135) <= layer1_outputs(8055);
    layer2_outputs(6136) <= layer1_outputs(1454);
    layer2_outputs(6137) <= (layer1_outputs(1968)) and not (layer1_outputs(9259));
    layer2_outputs(6138) <= not(layer1_outputs(198));
    layer2_outputs(6139) <= not(layer1_outputs(6200)) or (layer1_outputs(7584));
    layer2_outputs(6140) <= layer1_outputs(9200);
    layer2_outputs(6141) <= (layer1_outputs(8039)) xor (layer1_outputs(3507));
    layer2_outputs(6142) <= (layer1_outputs(3213)) xor (layer1_outputs(2994));
    layer2_outputs(6143) <= (layer1_outputs(8053)) and (layer1_outputs(7596));
    layer2_outputs(6144) <= (layer1_outputs(3485)) and not (layer1_outputs(1304));
    layer2_outputs(6145) <= layer1_outputs(5715);
    layer2_outputs(6146) <= layer1_outputs(2410);
    layer2_outputs(6147) <= not((layer1_outputs(836)) or (layer1_outputs(7026)));
    layer2_outputs(6148) <= not(layer1_outputs(3421));
    layer2_outputs(6149) <= not(layer1_outputs(7881)) or (layer1_outputs(1221));
    layer2_outputs(6150) <= layer1_outputs(3930);
    layer2_outputs(6151) <= not(layer1_outputs(1791));
    layer2_outputs(6152) <= not(layer1_outputs(4851));
    layer2_outputs(6153) <= not(layer1_outputs(2438));
    layer2_outputs(6154) <= not(layer1_outputs(8261));
    layer2_outputs(6155) <= not((layer1_outputs(4768)) and (layer1_outputs(5401)));
    layer2_outputs(6156) <= not(layer1_outputs(9812)) or (layer1_outputs(3948));
    layer2_outputs(6157) <= (layer1_outputs(10012)) and (layer1_outputs(7235));
    layer2_outputs(6158) <= layer1_outputs(92);
    layer2_outputs(6159) <= not(layer1_outputs(6537));
    layer2_outputs(6160) <= not(layer1_outputs(2874));
    layer2_outputs(6161) <= layer1_outputs(1589);
    layer2_outputs(6162) <= not(layer1_outputs(119));
    layer2_outputs(6163) <= (layer1_outputs(9287)) and (layer1_outputs(6759));
    layer2_outputs(6164) <= (layer1_outputs(7975)) and not (layer1_outputs(8728));
    layer2_outputs(6165) <= not(layer1_outputs(3985)) or (layer1_outputs(4976));
    layer2_outputs(6166) <= (layer1_outputs(4444)) and not (layer1_outputs(5873));
    layer2_outputs(6167) <= (layer1_outputs(7094)) and (layer1_outputs(8690));
    layer2_outputs(6168) <= (layer1_outputs(1827)) and not (layer1_outputs(8635));
    layer2_outputs(6169) <= (layer1_outputs(2136)) xor (layer1_outputs(9153));
    layer2_outputs(6170) <= not(layer1_outputs(3848)) or (layer1_outputs(1650));
    layer2_outputs(6171) <= not((layer1_outputs(4361)) and (layer1_outputs(1620)));
    layer2_outputs(6172) <= layer1_outputs(9666);
    layer2_outputs(6173) <= (layer1_outputs(8514)) and not (layer1_outputs(607));
    layer2_outputs(6174) <= not(layer1_outputs(2477));
    layer2_outputs(6175) <= not((layer1_outputs(6566)) xor (layer1_outputs(5617)));
    layer2_outputs(6176) <= layer1_outputs(1609);
    layer2_outputs(6177) <= not((layer1_outputs(1887)) xor (layer1_outputs(724)));
    layer2_outputs(6178) <= not(layer1_outputs(9966));
    layer2_outputs(6179) <= (layer1_outputs(3014)) xor (layer1_outputs(4066));
    layer2_outputs(6180) <= not((layer1_outputs(3779)) xor (layer1_outputs(4234)));
    layer2_outputs(6181) <= (layer1_outputs(6615)) and not (layer1_outputs(196));
    layer2_outputs(6182) <= not((layer1_outputs(2558)) xor (layer1_outputs(5778)));
    layer2_outputs(6183) <= (layer1_outputs(4690)) xor (layer1_outputs(1159));
    layer2_outputs(6184) <= not((layer1_outputs(5625)) and (layer1_outputs(1801)));
    layer2_outputs(6185) <= layer1_outputs(9124);
    layer2_outputs(6186) <= not((layer1_outputs(3765)) xor (layer1_outputs(9572)));
    layer2_outputs(6187) <= not(layer1_outputs(8302));
    layer2_outputs(6188) <= not(layer1_outputs(8120));
    layer2_outputs(6189) <= (layer1_outputs(6477)) and not (layer1_outputs(2872));
    layer2_outputs(6190) <= (layer1_outputs(7865)) and (layer1_outputs(4436));
    layer2_outputs(6191) <= layer1_outputs(1678);
    layer2_outputs(6192) <= not(layer1_outputs(9581));
    layer2_outputs(6193) <= not(layer1_outputs(5078)) or (layer1_outputs(4815));
    layer2_outputs(6194) <= (layer1_outputs(2258)) and (layer1_outputs(8717));
    layer2_outputs(6195) <= layer1_outputs(7);
    layer2_outputs(6196) <= not((layer1_outputs(6704)) or (layer1_outputs(3523)));
    layer2_outputs(6197) <= not(layer1_outputs(3444)) or (layer1_outputs(4681));
    layer2_outputs(6198) <= layer1_outputs(3320);
    layer2_outputs(6199) <= layer1_outputs(3816);
    layer2_outputs(6200) <= layer1_outputs(3782);
    layer2_outputs(6201) <= (layer1_outputs(2435)) and not (layer1_outputs(3363));
    layer2_outputs(6202) <= layer1_outputs(546);
    layer2_outputs(6203) <= (layer1_outputs(6770)) or (layer1_outputs(4507));
    layer2_outputs(6204) <= layer1_outputs(2094);
    layer2_outputs(6205) <= not((layer1_outputs(9706)) xor (layer1_outputs(7454)));
    layer2_outputs(6206) <= (layer1_outputs(1717)) or (layer1_outputs(7778));
    layer2_outputs(6207) <= not(layer1_outputs(9320));
    layer2_outputs(6208) <= layer1_outputs(7038);
    layer2_outputs(6209) <= layer1_outputs(7870);
    layer2_outputs(6210) <= not((layer1_outputs(943)) and (layer1_outputs(5193)));
    layer2_outputs(6211) <= (layer1_outputs(5836)) or (layer1_outputs(8374));
    layer2_outputs(6212) <= (layer1_outputs(1797)) xor (layer1_outputs(3445));
    layer2_outputs(6213) <= layer1_outputs(1608);
    layer2_outputs(6214) <= layer1_outputs(5520);
    layer2_outputs(6215) <= layer1_outputs(4327);
    layer2_outputs(6216) <= (layer1_outputs(50)) or (layer1_outputs(3450));
    layer2_outputs(6217) <= not(layer1_outputs(6));
    layer2_outputs(6218) <= not(layer1_outputs(567));
    layer2_outputs(6219) <= (layer1_outputs(7671)) and not (layer1_outputs(4275));
    layer2_outputs(6220) <= '1';
    layer2_outputs(6221) <= not(layer1_outputs(1997));
    layer2_outputs(6222) <= not(layer1_outputs(8377));
    layer2_outputs(6223) <= not(layer1_outputs(3757));
    layer2_outputs(6224) <= (layer1_outputs(8913)) and (layer1_outputs(1754));
    layer2_outputs(6225) <= not(layer1_outputs(6724)) or (layer1_outputs(10008));
    layer2_outputs(6226) <= layer1_outputs(825);
    layer2_outputs(6227) <= not((layer1_outputs(6880)) xor (layer1_outputs(9027)));
    layer2_outputs(6228) <= not(layer1_outputs(6377));
    layer2_outputs(6229) <= not(layer1_outputs(929));
    layer2_outputs(6230) <= layer1_outputs(8656);
    layer2_outputs(6231) <= not(layer1_outputs(8796));
    layer2_outputs(6232) <= not(layer1_outputs(91));
    layer2_outputs(6233) <= not((layer1_outputs(6210)) xor (layer1_outputs(6999)));
    layer2_outputs(6234) <= not(layer1_outputs(6541));
    layer2_outputs(6235) <= not(layer1_outputs(7718));
    layer2_outputs(6236) <= not((layer1_outputs(6247)) xor (layer1_outputs(442)));
    layer2_outputs(6237) <= (layer1_outputs(2657)) and (layer1_outputs(5365));
    layer2_outputs(6238) <= layer1_outputs(4884);
    layer2_outputs(6239) <= layer1_outputs(7200);
    layer2_outputs(6240) <= layer1_outputs(1854);
    layer2_outputs(6241) <= layer1_outputs(1502);
    layer2_outputs(6242) <= not(layer1_outputs(7852));
    layer2_outputs(6243) <= not(layer1_outputs(68)) or (layer1_outputs(59));
    layer2_outputs(6244) <= layer1_outputs(2191);
    layer2_outputs(6245) <= (layer1_outputs(1513)) xor (layer1_outputs(7045));
    layer2_outputs(6246) <= (layer1_outputs(7416)) and not (layer1_outputs(4980));
    layer2_outputs(6247) <= not((layer1_outputs(10140)) xor (layer1_outputs(7232)));
    layer2_outputs(6248) <= not(layer1_outputs(1538)) or (layer1_outputs(7257));
    layer2_outputs(6249) <= not(layer1_outputs(3677));
    layer2_outputs(6250) <= layer1_outputs(6918);
    layer2_outputs(6251) <= not((layer1_outputs(2284)) xor (layer1_outputs(1777)));
    layer2_outputs(6252) <= not(layer1_outputs(6191));
    layer2_outputs(6253) <= not(layer1_outputs(3360)) or (layer1_outputs(5));
    layer2_outputs(6254) <= (layer1_outputs(3053)) and not (layer1_outputs(5504));
    layer2_outputs(6255) <= not((layer1_outputs(7148)) and (layer1_outputs(5543)));
    layer2_outputs(6256) <= (layer1_outputs(9844)) xor (layer1_outputs(1923));
    layer2_outputs(6257) <= (layer1_outputs(2563)) and not (layer1_outputs(7676));
    layer2_outputs(6258) <= not(layer1_outputs(5665)) or (layer1_outputs(8487));
    layer2_outputs(6259) <= layer1_outputs(3579);
    layer2_outputs(6260) <= layer1_outputs(8169);
    layer2_outputs(6261) <= not(layer1_outputs(8821));
    layer2_outputs(6262) <= not(layer1_outputs(8400));
    layer2_outputs(6263) <= (layer1_outputs(7355)) and not (layer1_outputs(3836));
    layer2_outputs(6264) <= not(layer1_outputs(6243));
    layer2_outputs(6265) <= not((layer1_outputs(3342)) xor (layer1_outputs(562)));
    layer2_outputs(6266) <= not((layer1_outputs(3749)) and (layer1_outputs(4785)));
    layer2_outputs(6267) <= (layer1_outputs(1630)) and not (layer1_outputs(5060));
    layer2_outputs(6268) <= '0';
    layer2_outputs(6269) <= not((layer1_outputs(1660)) and (layer1_outputs(757)));
    layer2_outputs(6270) <= layer1_outputs(7508);
    layer2_outputs(6271) <= (layer1_outputs(8796)) xor (layer1_outputs(10081));
    layer2_outputs(6272) <= layer1_outputs(221);
    layer2_outputs(6273) <= not(layer1_outputs(497)) or (layer1_outputs(7922));
    layer2_outputs(6274) <= (layer1_outputs(2319)) and not (layer1_outputs(3835));
    layer2_outputs(6275) <= (layer1_outputs(4720)) and not (layer1_outputs(2488));
    layer2_outputs(6276) <= not(layer1_outputs(7000));
    layer2_outputs(6277) <= not(layer1_outputs(5394));
    layer2_outputs(6278) <= not(layer1_outputs(8907));
    layer2_outputs(6279) <= not(layer1_outputs(8604));
    layer2_outputs(6280) <= not(layer1_outputs(6953));
    layer2_outputs(6281) <= (layer1_outputs(4229)) and not (layer1_outputs(2143));
    layer2_outputs(6282) <= not((layer1_outputs(9231)) and (layer1_outputs(3832)));
    layer2_outputs(6283) <= (layer1_outputs(5122)) and (layer1_outputs(6168));
    layer2_outputs(6284) <= layer1_outputs(5708);
    layer2_outputs(6285) <= not((layer1_outputs(7742)) xor (layer1_outputs(6438)));
    layer2_outputs(6286) <= not(layer1_outputs(9667));
    layer2_outputs(6287) <= not(layer1_outputs(7317));
    layer2_outputs(6288) <= layer1_outputs(446);
    layer2_outputs(6289) <= layer1_outputs(3122);
    layer2_outputs(6290) <= not((layer1_outputs(7431)) xor (layer1_outputs(363)));
    layer2_outputs(6291) <= (layer1_outputs(2361)) and not (layer1_outputs(2475));
    layer2_outputs(6292) <= layer1_outputs(8229);
    layer2_outputs(6293) <= (layer1_outputs(9324)) xor (layer1_outputs(49));
    layer2_outputs(6294) <= not(layer1_outputs(8945));
    layer2_outputs(6295) <= layer1_outputs(5693);
    layer2_outputs(6296) <= not(layer1_outputs(5921));
    layer2_outputs(6297) <= not(layer1_outputs(3736));
    layer2_outputs(6298) <= not((layer1_outputs(4882)) or (layer1_outputs(4300)));
    layer2_outputs(6299) <= not((layer1_outputs(5216)) xor (layer1_outputs(5123)));
    layer2_outputs(6300) <= (layer1_outputs(10186)) xor (layer1_outputs(2758));
    layer2_outputs(6301) <= not((layer1_outputs(9367)) xor (layer1_outputs(2093)));
    layer2_outputs(6302) <= (layer1_outputs(3605)) and not (layer1_outputs(7019));
    layer2_outputs(6303) <= layer1_outputs(591);
    layer2_outputs(6304) <= layer1_outputs(9645);
    layer2_outputs(6305) <= not((layer1_outputs(4187)) xor (layer1_outputs(8502)));
    layer2_outputs(6306) <= not(layer1_outputs(822));
    layer2_outputs(6307) <= layer1_outputs(4492);
    layer2_outputs(6308) <= not((layer1_outputs(9746)) xor (layer1_outputs(4125)));
    layer2_outputs(6309) <= not(layer1_outputs(7939));
    layer2_outputs(6310) <= not(layer1_outputs(9640)) or (layer1_outputs(5282));
    layer2_outputs(6311) <= layer1_outputs(10185);
    layer2_outputs(6312) <= (layer1_outputs(708)) xor (layer1_outputs(5156));
    layer2_outputs(6313) <= not(layer1_outputs(8168)) or (layer1_outputs(761));
    layer2_outputs(6314) <= not(layer1_outputs(1014));
    layer2_outputs(6315) <= not((layer1_outputs(7777)) and (layer1_outputs(6238)));
    layer2_outputs(6316) <= (layer1_outputs(6633)) and not (layer1_outputs(1040));
    layer2_outputs(6317) <= layer1_outputs(1196);
    layer2_outputs(6318) <= not(layer1_outputs(3528)) or (layer1_outputs(7338));
    layer2_outputs(6319) <= not((layer1_outputs(1802)) or (layer1_outputs(8383)));
    layer2_outputs(6320) <= layer1_outputs(6209);
    layer2_outputs(6321) <= not(layer1_outputs(6923));
    layer2_outputs(6322) <= (layer1_outputs(4651)) and not (layer1_outputs(6403));
    layer2_outputs(6323) <= not(layer1_outputs(9033));
    layer2_outputs(6324) <= not(layer1_outputs(3089));
    layer2_outputs(6325) <= layer1_outputs(4939);
    layer2_outputs(6326) <= not((layer1_outputs(4815)) xor (layer1_outputs(5700)));
    layer2_outputs(6327) <= not(layer1_outputs(1)) or (layer1_outputs(1719));
    layer2_outputs(6328) <= (layer1_outputs(8388)) or (layer1_outputs(7881));
    layer2_outputs(6329) <= (layer1_outputs(604)) and not (layer1_outputs(3351));
    layer2_outputs(6330) <= layer1_outputs(4979);
    layer2_outputs(6331) <= layer1_outputs(1929);
    layer2_outputs(6332) <= layer1_outputs(2846);
    layer2_outputs(6333) <= not(layer1_outputs(4478));
    layer2_outputs(6334) <= not(layer1_outputs(1311));
    layer2_outputs(6335) <= (layer1_outputs(2436)) and not (layer1_outputs(2950));
    layer2_outputs(6336) <= not((layer1_outputs(6160)) xor (layer1_outputs(1745)));
    layer2_outputs(6337) <= layer1_outputs(9093);
    layer2_outputs(6338) <= (layer1_outputs(8521)) and (layer1_outputs(5229));
    layer2_outputs(6339) <= (layer1_outputs(7406)) or (layer1_outputs(7885));
    layer2_outputs(6340) <= not((layer1_outputs(536)) or (layer1_outputs(6831)));
    layer2_outputs(6341) <= not(layer1_outputs(6548));
    layer2_outputs(6342) <= layer1_outputs(765);
    layer2_outputs(6343) <= not((layer1_outputs(9169)) and (layer1_outputs(8652)));
    layer2_outputs(6344) <= layer1_outputs(286);
    layer2_outputs(6345) <= not(layer1_outputs(9293));
    layer2_outputs(6346) <= not(layer1_outputs(8167));
    layer2_outputs(6347) <= not(layer1_outputs(9934)) or (layer1_outputs(5577));
    layer2_outputs(6348) <= layer1_outputs(8914);
    layer2_outputs(6349) <= not(layer1_outputs(8791));
    layer2_outputs(6350) <= not(layer1_outputs(5908));
    layer2_outputs(6351) <= layer1_outputs(4440);
    layer2_outputs(6352) <= not((layer1_outputs(804)) xor (layer1_outputs(4524)));
    layer2_outputs(6353) <= not(layer1_outputs(4189));
    layer2_outputs(6354) <= not(layer1_outputs(256));
    layer2_outputs(6355) <= (layer1_outputs(746)) and (layer1_outputs(7271));
    layer2_outputs(6356) <= layer1_outputs(4667);
    layer2_outputs(6357) <= not(layer1_outputs(3));
    layer2_outputs(6358) <= not((layer1_outputs(3401)) or (layer1_outputs(1121)));
    layer2_outputs(6359) <= not(layer1_outputs(7943));
    layer2_outputs(6360) <= not((layer1_outputs(4578)) and (layer1_outputs(9091)));
    layer2_outputs(6361) <= (layer1_outputs(5457)) xor (layer1_outputs(4421));
    layer2_outputs(6362) <= layer1_outputs(2302);
    layer2_outputs(6363) <= layer1_outputs(7665);
    layer2_outputs(6364) <= not(layer1_outputs(5474));
    layer2_outputs(6365) <= not((layer1_outputs(63)) or (layer1_outputs(156)));
    layer2_outputs(6366) <= layer1_outputs(9063);
    layer2_outputs(6367) <= (layer1_outputs(9768)) or (layer1_outputs(8531));
    layer2_outputs(6368) <= not(layer1_outputs(2862)) or (layer1_outputs(3233));
    layer2_outputs(6369) <= not(layer1_outputs(6914));
    layer2_outputs(6370) <= '1';
    layer2_outputs(6371) <= layer1_outputs(5083);
    layer2_outputs(6372) <= '1';
    layer2_outputs(6373) <= not(layer1_outputs(4876));
    layer2_outputs(6374) <= layer1_outputs(3857);
    layer2_outputs(6375) <= '0';
    layer2_outputs(6376) <= not(layer1_outputs(4710));
    layer2_outputs(6377) <= not(layer1_outputs(9078));
    layer2_outputs(6378) <= not(layer1_outputs(8271));
    layer2_outputs(6379) <= not(layer1_outputs(8992)) or (layer1_outputs(10003));
    layer2_outputs(6380) <= layer1_outputs(6366);
    layer2_outputs(6381) <= not((layer1_outputs(1662)) or (layer1_outputs(9872)));
    layer2_outputs(6382) <= not(layer1_outputs(1345));
    layer2_outputs(6383) <= not(layer1_outputs(9753));
    layer2_outputs(6384) <= not((layer1_outputs(6955)) xor (layer1_outputs(1032)));
    layer2_outputs(6385) <= (layer1_outputs(9658)) xor (layer1_outputs(1659));
    layer2_outputs(6386) <= not((layer1_outputs(5889)) xor (layer1_outputs(3237)));
    layer2_outputs(6387) <= layer1_outputs(5259);
    layer2_outputs(6388) <= not(layer1_outputs(407));
    layer2_outputs(6389) <= layer1_outputs(1746);
    layer2_outputs(6390) <= not(layer1_outputs(4018));
    layer2_outputs(6391) <= layer1_outputs(8520);
    layer2_outputs(6392) <= layer1_outputs(6841);
    layer2_outputs(6393) <= (layer1_outputs(9874)) and (layer1_outputs(1232));
    layer2_outputs(6394) <= not((layer1_outputs(6144)) xor (layer1_outputs(4245)));
    layer2_outputs(6395) <= (layer1_outputs(733)) and not (layer1_outputs(9823));
    layer2_outputs(6396) <= layer1_outputs(5302);
    layer2_outputs(6397) <= (layer1_outputs(4895)) and not (layer1_outputs(4765));
    layer2_outputs(6398) <= not(layer1_outputs(5663));
    layer2_outputs(6399) <= not(layer1_outputs(9406));
    layer2_outputs(6400) <= (layer1_outputs(10219)) xor (layer1_outputs(5688));
    layer2_outputs(6401) <= '0';
    layer2_outputs(6402) <= not(layer1_outputs(6331));
    layer2_outputs(6403) <= not(layer1_outputs(1775));
    layer2_outputs(6404) <= not((layer1_outputs(4661)) xor (layer1_outputs(2009)));
    layer2_outputs(6405) <= not(layer1_outputs(10175));
    layer2_outputs(6406) <= (layer1_outputs(252)) and not (layer1_outputs(9251));
    layer2_outputs(6407) <= (layer1_outputs(9990)) or (layer1_outputs(8946));
    layer2_outputs(6408) <= (layer1_outputs(6915)) and not (layer1_outputs(9434));
    layer2_outputs(6409) <= not(layer1_outputs(1956));
    layer2_outputs(6410) <= not(layer1_outputs(7329)) or (layer1_outputs(6325));
    layer2_outputs(6411) <= layer1_outputs(10196);
    layer2_outputs(6412) <= (layer1_outputs(103)) xor (layer1_outputs(9945));
    layer2_outputs(6413) <= (layer1_outputs(3310)) and not (layer1_outputs(3681));
    layer2_outputs(6414) <= (layer1_outputs(5930)) and (layer1_outputs(8424));
    layer2_outputs(6415) <= not((layer1_outputs(915)) and (layer1_outputs(10097)));
    layer2_outputs(6416) <= (layer1_outputs(4111)) and (layer1_outputs(1201));
    layer2_outputs(6417) <= not(layer1_outputs(8138));
    layer2_outputs(6418) <= not(layer1_outputs(177));
    layer2_outputs(6419) <= not(layer1_outputs(7366));
    layer2_outputs(6420) <= not((layer1_outputs(4212)) xor (layer1_outputs(563)));
    layer2_outputs(6421) <= layer1_outputs(1775);
    layer2_outputs(6422) <= not(layer1_outputs(5473)) or (layer1_outputs(5944));
    layer2_outputs(6423) <= not((layer1_outputs(9646)) and (layer1_outputs(4228)));
    layer2_outputs(6424) <= not(layer1_outputs(6590));
    layer2_outputs(6425) <= (layer1_outputs(9549)) and not (layer1_outputs(9325));
    layer2_outputs(6426) <= not(layer1_outputs(5319));
    layer2_outputs(6427) <= not((layer1_outputs(9837)) or (layer1_outputs(5344)));
    layer2_outputs(6428) <= not(layer1_outputs(3570));
    layer2_outputs(6429) <= not(layer1_outputs(2949));
    layer2_outputs(6430) <= layer1_outputs(7450);
    layer2_outputs(6431) <= not(layer1_outputs(3090)) or (layer1_outputs(5864));
    layer2_outputs(6432) <= not(layer1_outputs(5988));
    layer2_outputs(6433) <= not(layer1_outputs(2867));
    layer2_outputs(6434) <= not((layer1_outputs(376)) xor (layer1_outputs(6654)));
    layer2_outputs(6435) <= layer1_outputs(141);
    layer2_outputs(6436) <= not(layer1_outputs(451)) or (layer1_outputs(7163));
    layer2_outputs(6437) <= (layer1_outputs(7578)) or (layer1_outputs(9186));
    layer2_outputs(6438) <= layer1_outputs(4365);
    layer2_outputs(6439) <= layer1_outputs(7127);
    layer2_outputs(6440) <= (layer1_outputs(781)) xor (layer1_outputs(7422));
    layer2_outputs(6441) <= (layer1_outputs(6408)) or (layer1_outputs(1423));
    layer2_outputs(6442) <= not(layer1_outputs(2159));
    layer2_outputs(6443) <= not((layer1_outputs(879)) and (layer1_outputs(8860)));
    layer2_outputs(6444) <= not(layer1_outputs(8159));
    layer2_outputs(6445) <= layer1_outputs(5253);
    layer2_outputs(6446) <= (layer1_outputs(3136)) and not (layer1_outputs(9376));
    layer2_outputs(6447) <= not(layer1_outputs(5776));
    layer2_outputs(6448) <= (layer1_outputs(8140)) and (layer1_outputs(8526));
    layer2_outputs(6449) <= not(layer1_outputs(8550));
    layer2_outputs(6450) <= not((layer1_outputs(1447)) xor (layer1_outputs(5878)));
    layer2_outputs(6451) <= (layer1_outputs(4746)) and (layer1_outputs(1149));
    layer2_outputs(6452) <= not(layer1_outputs(900));
    layer2_outputs(6453) <= layer1_outputs(6916);
    layer2_outputs(6454) <= layer1_outputs(7650);
    layer2_outputs(6455) <= not(layer1_outputs(9451));
    layer2_outputs(6456) <= not(layer1_outputs(1633));
    layer2_outputs(6457) <= not(layer1_outputs(3968));
    layer2_outputs(6458) <= not((layer1_outputs(9558)) and (layer1_outputs(5763)));
    layer2_outputs(6459) <= not((layer1_outputs(190)) xor (layer1_outputs(6488)));
    layer2_outputs(6460) <= layer1_outputs(9834);
    layer2_outputs(6461) <= not(layer1_outputs(9510));
    layer2_outputs(6462) <= (layer1_outputs(7077)) and not (layer1_outputs(4638));
    layer2_outputs(6463) <= (layer1_outputs(2930)) and not (layer1_outputs(6703));
    layer2_outputs(6464) <= not(layer1_outputs(2129));
    layer2_outputs(6465) <= layer1_outputs(3006);
    layer2_outputs(6466) <= not(layer1_outputs(3163));
    layer2_outputs(6467) <= not(layer1_outputs(7529));
    layer2_outputs(6468) <= (layer1_outputs(4899)) or (layer1_outputs(10174));
    layer2_outputs(6469) <= not((layer1_outputs(8751)) or (layer1_outputs(1514)));
    layer2_outputs(6470) <= not((layer1_outputs(1499)) xor (layer1_outputs(6256)));
    layer2_outputs(6471) <= layer1_outputs(8222);
    layer2_outputs(6472) <= not((layer1_outputs(8236)) and (layer1_outputs(5546)));
    layer2_outputs(6473) <= (layer1_outputs(3512)) and not (layer1_outputs(3204));
    layer2_outputs(6474) <= not((layer1_outputs(597)) xor (layer1_outputs(5175)));
    layer2_outputs(6475) <= (layer1_outputs(8766)) and not (layer1_outputs(5265));
    layer2_outputs(6476) <= layer1_outputs(8339);
    layer2_outputs(6477) <= (layer1_outputs(10084)) and not (layer1_outputs(5016));
    layer2_outputs(6478) <= layer1_outputs(8881);
    layer2_outputs(6479) <= not(layer1_outputs(839)) or (layer1_outputs(2977));
    layer2_outputs(6480) <= layer1_outputs(1986);
    layer2_outputs(6481) <= not(layer1_outputs(2651));
    layer2_outputs(6482) <= not(layer1_outputs(1832));
    layer2_outputs(6483) <= layer1_outputs(3124);
    layer2_outputs(6484) <= (layer1_outputs(6244)) xor (layer1_outputs(8406));
    layer2_outputs(6485) <= (layer1_outputs(5133)) or (layer1_outputs(951));
    layer2_outputs(6486) <= not((layer1_outputs(10160)) xor (layer1_outputs(9560)));
    layer2_outputs(6487) <= not((layer1_outputs(4944)) or (layer1_outputs(1275)));
    layer2_outputs(6488) <= not((layer1_outputs(903)) or (layer1_outputs(1054)));
    layer2_outputs(6489) <= (layer1_outputs(3676)) and not (layer1_outputs(891));
    layer2_outputs(6490) <= (layer1_outputs(9550)) xor (layer1_outputs(6538));
    layer2_outputs(6491) <= '1';
    layer2_outputs(6492) <= layer1_outputs(9884);
    layer2_outputs(6493) <= layer1_outputs(2074);
    layer2_outputs(6494) <= (layer1_outputs(3510)) and not (layer1_outputs(3321));
    layer2_outputs(6495) <= layer1_outputs(2587);
    layer2_outputs(6496) <= layer1_outputs(341);
    layer2_outputs(6497) <= (layer1_outputs(9385)) and not (layer1_outputs(10043));
    layer2_outputs(6498) <= not((layer1_outputs(445)) and (layer1_outputs(8019)));
    layer2_outputs(6499) <= not((layer1_outputs(7594)) and (layer1_outputs(714)));
    layer2_outputs(6500) <= (layer1_outputs(1610)) and not (layer1_outputs(6598));
    layer2_outputs(6501) <= not(layer1_outputs(6358)) or (layer1_outputs(4549));
    layer2_outputs(6502) <= (layer1_outputs(327)) and not (layer1_outputs(4802));
    layer2_outputs(6503) <= (layer1_outputs(2708)) and not (layer1_outputs(267));
    layer2_outputs(6504) <= not(layer1_outputs(501));
    layer2_outputs(6505) <= not(layer1_outputs(7615));
    layer2_outputs(6506) <= (layer1_outputs(2027)) and not (layer1_outputs(7483));
    layer2_outputs(6507) <= not((layer1_outputs(9558)) and (layer1_outputs(42)));
    layer2_outputs(6508) <= layer1_outputs(3902);
    layer2_outputs(6509) <= (layer1_outputs(9489)) and not (layer1_outputs(5067));
    layer2_outputs(6510) <= layer1_outputs(5971);
    layer2_outputs(6511) <= (layer1_outputs(8271)) and not (layer1_outputs(3171));
    layer2_outputs(6512) <= (layer1_outputs(4700)) and (layer1_outputs(2374));
    layer2_outputs(6513) <= layer1_outputs(4237);
    layer2_outputs(6514) <= (layer1_outputs(791)) xor (layer1_outputs(10070));
    layer2_outputs(6515) <= not(layer1_outputs(5403));
    layer2_outputs(6516) <= not((layer1_outputs(419)) or (layer1_outputs(2826)));
    layer2_outputs(6517) <= (layer1_outputs(1344)) or (layer1_outputs(9207));
    layer2_outputs(6518) <= not((layer1_outputs(1769)) and (layer1_outputs(7045)));
    layer2_outputs(6519) <= not(layer1_outputs(203));
    layer2_outputs(6520) <= (layer1_outputs(656)) xor (layer1_outputs(6211));
    layer2_outputs(6521) <= '0';
    layer2_outputs(6522) <= (layer1_outputs(4831)) xor (layer1_outputs(8823));
    layer2_outputs(6523) <= layer1_outputs(577);
    layer2_outputs(6524) <= (layer1_outputs(3007)) and not (layer1_outputs(9593));
    layer2_outputs(6525) <= not((layer1_outputs(8350)) xor (layer1_outputs(460)));
    layer2_outputs(6526) <= layer1_outputs(7988);
    layer2_outputs(6527) <= not(layer1_outputs(4735));
    layer2_outputs(6528) <= (layer1_outputs(9981)) or (layer1_outputs(4571));
    layer2_outputs(6529) <= not(layer1_outputs(9591));
    layer2_outputs(6530) <= (layer1_outputs(3631)) and not (layer1_outputs(6245));
    layer2_outputs(6531) <= not(layer1_outputs(9125));
    layer2_outputs(6532) <= (layer1_outputs(4913)) and (layer1_outputs(9142));
    layer2_outputs(6533) <= (layer1_outputs(1886)) and not (layer1_outputs(6559));
    layer2_outputs(6534) <= layer1_outputs(614);
    layer2_outputs(6535) <= layer1_outputs(9134);
    layer2_outputs(6536) <= (layer1_outputs(3700)) or (layer1_outputs(8575));
    layer2_outputs(6537) <= (layer1_outputs(5513)) xor (layer1_outputs(6638));
    layer2_outputs(6538) <= (layer1_outputs(730)) and not (layer1_outputs(663));
    layer2_outputs(6539) <= (layer1_outputs(10025)) xor (layer1_outputs(6021));
    layer2_outputs(6540) <= (layer1_outputs(5787)) and not (layer1_outputs(9887));
    layer2_outputs(6541) <= (layer1_outputs(9468)) and (layer1_outputs(9480));
    layer2_outputs(6542) <= not(layer1_outputs(5361));
    layer2_outputs(6543) <= not((layer1_outputs(4662)) or (layer1_outputs(6192)));
    layer2_outputs(6544) <= layer1_outputs(3186);
    layer2_outputs(6545) <= not(layer1_outputs(1022));
    layer2_outputs(6546) <= not(layer1_outputs(162));
    layer2_outputs(6547) <= not((layer1_outputs(5564)) and (layer1_outputs(4838)));
    layer2_outputs(6548) <= not(layer1_outputs(4399));
    layer2_outputs(6549) <= (layer1_outputs(3374)) or (layer1_outputs(8864));
    layer2_outputs(6550) <= layer1_outputs(3740);
    layer2_outputs(6551) <= not(layer1_outputs(2449));
    layer2_outputs(6552) <= (layer1_outputs(1427)) and not (layer1_outputs(8181));
    layer2_outputs(6553) <= not(layer1_outputs(3806));
    layer2_outputs(6554) <= not(layer1_outputs(2541));
    layer2_outputs(6555) <= not((layer1_outputs(689)) and (layer1_outputs(9227)));
    layer2_outputs(6556) <= not(layer1_outputs(9670));
    layer2_outputs(6557) <= not(layer1_outputs(6149));
    layer2_outputs(6558) <= (layer1_outputs(9249)) and (layer1_outputs(7646));
    layer2_outputs(6559) <= not(layer1_outputs(2835)) or (layer1_outputs(2302));
    layer2_outputs(6560) <= not(layer1_outputs(8059));
    layer2_outputs(6561) <= layer1_outputs(2921);
    layer2_outputs(6562) <= layer1_outputs(8757);
    layer2_outputs(6563) <= not(layer1_outputs(605)) or (layer1_outputs(2386));
    layer2_outputs(6564) <= (layer1_outputs(8509)) and not (layer1_outputs(498));
    layer2_outputs(6565) <= layer1_outputs(5501);
    layer2_outputs(6566) <= layer1_outputs(715);
    layer2_outputs(6567) <= layer1_outputs(1722);
    layer2_outputs(6568) <= layer1_outputs(9748);
    layer2_outputs(6569) <= not(layer1_outputs(681));
    layer2_outputs(6570) <= not((layer1_outputs(7487)) or (layer1_outputs(7638)));
    layer2_outputs(6571) <= (layer1_outputs(9165)) xor (layer1_outputs(3860));
    layer2_outputs(6572) <= (layer1_outputs(10031)) and (layer1_outputs(9601));
    layer2_outputs(6573) <= layer1_outputs(5365);
    layer2_outputs(6574) <= (layer1_outputs(2609)) or (layer1_outputs(3387));
    layer2_outputs(6575) <= layer1_outputs(4890);
    layer2_outputs(6576) <= not(layer1_outputs(2879));
    layer2_outputs(6577) <= not(layer1_outputs(7273)) or (layer1_outputs(4983));
    layer2_outputs(6578) <= (layer1_outputs(8843)) and not (layer1_outputs(5187));
    layer2_outputs(6579) <= not(layer1_outputs(2164));
    layer2_outputs(6580) <= not(layer1_outputs(5126)) or (layer1_outputs(2040));
    layer2_outputs(6581) <= not((layer1_outputs(8993)) xor (layer1_outputs(9985)));
    layer2_outputs(6582) <= layer1_outputs(9707);
    layer2_outputs(6583) <= not(layer1_outputs(208));
    layer2_outputs(6584) <= not(layer1_outputs(193)) or (layer1_outputs(7525));
    layer2_outputs(6585) <= (layer1_outputs(6293)) xor (layer1_outputs(9979));
    layer2_outputs(6586) <= layer1_outputs(8215);
    layer2_outputs(6587) <= (layer1_outputs(3655)) or (layer1_outputs(262));
    layer2_outputs(6588) <= layer1_outputs(2149);
    layer2_outputs(6589) <= not(layer1_outputs(3430));
    layer2_outputs(6590) <= not((layer1_outputs(569)) and (layer1_outputs(2208)));
    layer2_outputs(6591) <= layer1_outputs(2984);
    layer2_outputs(6592) <= '0';
    layer2_outputs(6593) <= not(layer1_outputs(4643)) or (layer1_outputs(3628));
    layer2_outputs(6594) <= layer1_outputs(6350);
    layer2_outputs(6595) <= not(layer1_outputs(875));
    layer2_outputs(6596) <= layer1_outputs(8149);
    layer2_outputs(6597) <= not((layer1_outputs(8805)) and (layer1_outputs(3921)));
    layer2_outputs(6598) <= not(layer1_outputs(6741));
    layer2_outputs(6599) <= (layer1_outputs(2595)) and not (layer1_outputs(2508));
    layer2_outputs(6600) <= not((layer1_outputs(5378)) xor (layer1_outputs(175)));
    layer2_outputs(6601) <= not((layer1_outputs(8263)) or (layer1_outputs(5265)));
    layer2_outputs(6602) <= layer1_outputs(292);
    layer2_outputs(6603) <= layer1_outputs(5149);
    layer2_outputs(6604) <= not(layer1_outputs(4582));
    layer2_outputs(6605) <= not((layer1_outputs(4673)) and (layer1_outputs(4756)));
    layer2_outputs(6606) <= '1';
    layer2_outputs(6607) <= not((layer1_outputs(7806)) or (layer1_outputs(6297)));
    layer2_outputs(6608) <= layer1_outputs(60);
    layer2_outputs(6609) <= (layer1_outputs(9721)) and not (layer1_outputs(2082));
    layer2_outputs(6610) <= not(layer1_outputs(6649));
    layer2_outputs(6611) <= not(layer1_outputs(9351));
    layer2_outputs(6612) <= not(layer1_outputs(6939)) or (layer1_outputs(5998));
    layer2_outputs(6613) <= not(layer1_outputs(1880));
    layer2_outputs(6614) <= (layer1_outputs(5979)) xor (layer1_outputs(322));
    layer2_outputs(6615) <= not(layer1_outputs(6289)) or (layer1_outputs(5746));
    layer2_outputs(6616) <= (layer1_outputs(1328)) and not (layer1_outputs(7827));
    layer2_outputs(6617) <= not(layer1_outputs(3265)) or (layer1_outputs(9543));
    layer2_outputs(6618) <= not(layer1_outputs(3423)) or (layer1_outputs(59));
    layer2_outputs(6619) <= not((layer1_outputs(8603)) or (layer1_outputs(6582)));
    layer2_outputs(6620) <= (layer1_outputs(5209)) or (layer1_outputs(5491));
    layer2_outputs(6621) <= not(layer1_outputs(280)) or (layer1_outputs(173));
    layer2_outputs(6622) <= not((layer1_outputs(7833)) or (layer1_outputs(4930)));
    layer2_outputs(6623) <= layer1_outputs(8599);
    layer2_outputs(6624) <= (layer1_outputs(2841)) and not (layer1_outputs(7470));
    layer2_outputs(6625) <= (layer1_outputs(9429)) and (layer1_outputs(5029));
    layer2_outputs(6626) <= (layer1_outputs(7358)) xor (layer1_outputs(748));
    layer2_outputs(6627) <= (layer1_outputs(10184)) xor (layer1_outputs(5430));
    layer2_outputs(6628) <= (layer1_outputs(2109)) and (layer1_outputs(687));
    layer2_outputs(6629) <= not(layer1_outputs(3669));
    layer2_outputs(6630) <= not(layer1_outputs(4416)) or (layer1_outputs(9578));
    layer2_outputs(6631) <= not((layer1_outputs(7877)) and (layer1_outputs(9805)));
    layer2_outputs(6632) <= (layer1_outputs(5372)) and not (layer1_outputs(2834));
    layer2_outputs(6633) <= layer1_outputs(9000);
    layer2_outputs(6634) <= layer1_outputs(1108);
    layer2_outputs(6635) <= not(layer1_outputs(3527)) or (layer1_outputs(5649));
    layer2_outputs(6636) <= not(layer1_outputs(3607));
    layer2_outputs(6637) <= not(layer1_outputs(7882));
    layer2_outputs(6638) <= (layer1_outputs(8543)) and not (layer1_outputs(2649));
    layer2_outputs(6639) <= layer1_outputs(9615);
    layer2_outputs(6640) <= (layer1_outputs(7911)) and not (layer1_outputs(1685));
    layer2_outputs(6641) <= not((layer1_outputs(31)) or (layer1_outputs(8163)));
    layer2_outputs(6642) <= (layer1_outputs(4686)) and (layer1_outputs(4842));
    layer2_outputs(6643) <= layer1_outputs(6922);
    layer2_outputs(6644) <= (layer1_outputs(8324)) and (layer1_outputs(3335));
    layer2_outputs(6645) <= not((layer1_outputs(3589)) xor (layer1_outputs(6732)));
    layer2_outputs(6646) <= not(layer1_outputs(7868));
    layer2_outputs(6647) <= layer1_outputs(218);
    layer2_outputs(6648) <= layer1_outputs(9330);
    layer2_outputs(6649) <= layer1_outputs(7946);
    layer2_outputs(6650) <= not(layer1_outputs(9629));
    layer2_outputs(6651) <= (layer1_outputs(3411)) or (layer1_outputs(10042));
    layer2_outputs(6652) <= (layer1_outputs(1874)) and not (layer1_outputs(5651));
    layer2_outputs(6653) <= not(layer1_outputs(8211)) or (layer1_outputs(3644));
    layer2_outputs(6654) <= layer1_outputs(685);
    layer2_outputs(6655) <= layer1_outputs(3582);
    layer2_outputs(6656) <= layer1_outputs(8137);
    layer2_outputs(6657) <= layer1_outputs(19);
    layer2_outputs(6658) <= layer1_outputs(3751);
    layer2_outputs(6659) <= not(layer1_outputs(3021));
    layer2_outputs(6660) <= not(layer1_outputs(2802));
    layer2_outputs(6661) <= layer1_outputs(4086);
    layer2_outputs(6662) <= not(layer1_outputs(35)) or (layer1_outputs(6102));
    layer2_outputs(6663) <= layer1_outputs(5954);
    layer2_outputs(6664) <= not(layer1_outputs(8997));
    layer2_outputs(6665) <= not(layer1_outputs(826));
    layer2_outputs(6666) <= not(layer1_outputs(5441));
    layer2_outputs(6667) <= not(layer1_outputs(9819)) or (layer1_outputs(1245));
    layer2_outputs(6668) <= not(layer1_outputs(9070));
    layer2_outputs(6669) <= layer1_outputs(1479);
    layer2_outputs(6670) <= layer1_outputs(5482);
    layer2_outputs(6671) <= (layer1_outputs(8093)) or (layer1_outputs(8105));
    layer2_outputs(6672) <= '0';
    layer2_outputs(6673) <= layer1_outputs(5972);
    layer2_outputs(6674) <= not(layer1_outputs(4976)) or (layer1_outputs(7723));
    layer2_outputs(6675) <= layer1_outputs(2112);
    layer2_outputs(6676) <= not(layer1_outputs(1212));
    layer2_outputs(6677) <= layer1_outputs(6622);
    layer2_outputs(6678) <= (layer1_outputs(5371)) and not (layer1_outputs(2165));
    layer2_outputs(6679) <= (layer1_outputs(3590)) and not (layer1_outputs(6917));
    layer2_outputs(6680) <= not(layer1_outputs(6196));
    layer2_outputs(6681) <= not(layer1_outputs(1200));
    layer2_outputs(6682) <= layer1_outputs(7549);
    layer2_outputs(6683) <= not(layer1_outputs(7167));
    layer2_outputs(6684) <= not(layer1_outputs(3283));
    layer2_outputs(6685) <= layer1_outputs(5785);
    layer2_outputs(6686) <= layer1_outputs(4344);
    layer2_outputs(6687) <= not(layer1_outputs(6333));
    layer2_outputs(6688) <= not(layer1_outputs(8485));
    layer2_outputs(6689) <= (layer1_outputs(2192)) and not (layer1_outputs(8368));
    layer2_outputs(6690) <= layer1_outputs(8867);
    layer2_outputs(6691) <= layer1_outputs(9002);
    layer2_outputs(6692) <= not(layer1_outputs(4182)) or (layer1_outputs(723));
    layer2_outputs(6693) <= not(layer1_outputs(3261)) or (layer1_outputs(6128));
    layer2_outputs(6694) <= not(layer1_outputs(3427)) or (layer1_outputs(7283));
    layer2_outputs(6695) <= not(layer1_outputs(3778));
    layer2_outputs(6696) <= not((layer1_outputs(6447)) and (layer1_outputs(7407)));
    layer2_outputs(6697) <= layer1_outputs(3164);
    layer2_outputs(6698) <= '0';
    layer2_outputs(6699) <= (layer1_outputs(1324)) or (layer1_outputs(1367));
    layer2_outputs(6700) <= not((layer1_outputs(9829)) or (layer1_outputs(275)));
    layer2_outputs(6701) <= layer1_outputs(8952);
    layer2_outputs(6702) <= (layer1_outputs(5646)) and not (layer1_outputs(388));
    layer2_outputs(6703) <= not(layer1_outputs(2476)) or (layer1_outputs(5443));
    layer2_outputs(6704) <= (layer1_outputs(6544)) xor (layer1_outputs(6920));
    layer2_outputs(6705) <= not(layer1_outputs(6491)) or (layer1_outputs(5419));
    layer2_outputs(6706) <= not(layer1_outputs(3037));
    layer2_outputs(6707) <= not((layer1_outputs(1877)) xor (layer1_outputs(633)));
    layer2_outputs(6708) <= (layer1_outputs(815)) and not (layer1_outputs(173));
    layer2_outputs(6709) <= layer1_outputs(3595);
    layer2_outputs(6710) <= layer1_outputs(2383);
    layer2_outputs(6711) <= not(layer1_outputs(8009));
    layer2_outputs(6712) <= layer1_outputs(1763);
    layer2_outputs(6713) <= (layer1_outputs(3188)) or (layer1_outputs(7687));
    layer2_outputs(6714) <= layer1_outputs(7905);
    layer2_outputs(6715) <= not(layer1_outputs(2659));
    layer2_outputs(6716) <= not(layer1_outputs(6271));
    layer2_outputs(6717) <= not(layer1_outputs(1435));
    layer2_outputs(6718) <= not(layer1_outputs(827)) or (layer1_outputs(6853));
    layer2_outputs(6719) <= not((layer1_outputs(9640)) or (layer1_outputs(456)));
    layer2_outputs(6720) <= layer1_outputs(10002);
    layer2_outputs(6721) <= not(layer1_outputs(7402));
    layer2_outputs(6722) <= layer1_outputs(9900);
    layer2_outputs(6723) <= not(layer1_outputs(5280)) or (layer1_outputs(1244));
    layer2_outputs(6724) <= (layer1_outputs(6885)) xor (layer1_outputs(8427));
    layer2_outputs(6725) <= not((layer1_outputs(7404)) or (layer1_outputs(546)));
    layer2_outputs(6726) <= not(layer1_outputs(2258));
    layer2_outputs(6727) <= not(layer1_outputs(1629));
    layer2_outputs(6728) <= (layer1_outputs(161)) and not (layer1_outputs(1913));
    layer2_outputs(6729) <= not(layer1_outputs(6961));
    layer2_outputs(6730) <= not(layer1_outputs(664));
    layer2_outputs(6731) <= (layer1_outputs(83)) or (layer1_outputs(8058));
    layer2_outputs(6732) <= not(layer1_outputs(1483)) or (layer1_outputs(7810));
    layer2_outputs(6733) <= layer1_outputs(3229);
    layer2_outputs(6734) <= layer1_outputs(4828);
    layer2_outputs(6735) <= layer1_outputs(1291);
    layer2_outputs(6736) <= layer1_outputs(6997);
    layer2_outputs(6737) <= not(layer1_outputs(10007));
    layer2_outputs(6738) <= layer1_outputs(772);
    layer2_outputs(6739) <= '0';
    layer2_outputs(6740) <= layer1_outputs(8321);
    layer2_outputs(6741) <= not(layer1_outputs(6309)) or (layer1_outputs(1041));
    layer2_outputs(6742) <= layer1_outputs(2031);
    layer2_outputs(6743) <= not(layer1_outputs(9717)) or (layer1_outputs(522));
    layer2_outputs(6744) <= (layer1_outputs(7227)) and not (layer1_outputs(516));
    layer2_outputs(6745) <= not((layer1_outputs(4613)) xor (layer1_outputs(1240)));
    layer2_outputs(6746) <= not(layer1_outputs(5669));
    layer2_outputs(6747) <= layer1_outputs(3474);
    layer2_outputs(6748) <= not(layer1_outputs(1241)) or (layer1_outputs(3437));
    layer2_outputs(6749) <= (layer1_outputs(7677)) and not (layer1_outputs(238));
    layer2_outputs(6750) <= (layer1_outputs(2621)) or (layer1_outputs(7493));
    layer2_outputs(6751) <= (layer1_outputs(8401)) and not (layer1_outputs(5702));
    layer2_outputs(6752) <= layer1_outputs(6874);
    layer2_outputs(6753) <= not(layer1_outputs(339));
    layer2_outputs(6754) <= (layer1_outputs(2207)) and (layer1_outputs(7903));
    layer2_outputs(6755) <= layer1_outputs(8673);
    layer2_outputs(6756) <= not((layer1_outputs(959)) or (layer1_outputs(2801)));
    layer2_outputs(6757) <= (layer1_outputs(3598)) and not (layer1_outputs(3842));
    layer2_outputs(6758) <= not(layer1_outputs(1233));
    layer2_outputs(6759) <= (layer1_outputs(4123)) and (layer1_outputs(843));
    layer2_outputs(6760) <= not(layer1_outputs(10083));
    layer2_outputs(6761) <= layer1_outputs(7693);
    layer2_outputs(6762) <= not((layer1_outputs(5880)) xor (layer1_outputs(7868)));
    layer2_outputs(6763) <= not((layer1_outputs(5186)) or (layer1_outputs(7751)));
    layer2_outputs(6764) <= (layer1_outputs(5529)) and not (layer1_outputs(8134));
    layer2_outputs(6765) <= (layer1_outputs(1757)) or (layer1_outputs(8064));
    layer2_outputs(6766) <= layer1_outputs(4160);
    layer2_outputs(6767) <= not(layer1_outputs(3334));
    layer2_outputs(6768) <= not((layer1_outputs(709)) xor (layer1_outputs(2611)));
    layer2_outputs(6769) <= (layer1_outputs(2298)) and (layer1_outputs(7144));
    layer2_outputs(6770) <= (layer1_outputs(6402)) xor (layer1_outputs(5569));
    layer2_outputs(6771) <= layer1_outputs(5785);
    layer2_outputs(6772) <= not((layer1_outputs(4113)) or (layer1_outputs(7870)));
    layer2_outputs(6773) <= not(layer1_outputs(5784));
    layer2_outputs(6774) <= (layer1_outputs(3370)) xor (layer1_outputs(1626));
    layer2_outputs(6775) <= not(layer1_outputs(8446));
    layer2_outputs(6776) <= (layer1_outputs(462)) xor (layer1_outputs(4101));
    layer2_outputs(6777) <= layer1_outputs(4457);
    layer2_outputs(6778) <= layer1_outputs(152);
    layer2_outputs(6779) <= layer1_outputs(6244);
    layer2_outputs(6780) <= (layer1_outputs(7552)) xor (layer1_outputs(8617));
    layer2_outputs(6781) <= not(layer1_outputs(9699));
    layer2_outputs(6782) <= not(layer1_outputs(3926));
    layer2_outputs(6783) <= not(layer1_outputs(382));
    layer2_outputs(6784) <= not((layer1_outputs(7628)) and (layer1_outputs(4935)));
    layer2_outputs(6785) <= not((layer1_outputs(987)) xor (layer1_outputs(4687)));
    layer2_outputs(6786) <= layer1_outputs(621);
    layer2_outputs(6787) <= (layer1_outputs(8351)) or (layer1_outputs(5093));
    layer2_outputs(6788) <= (layer1_outputs(3056)) xor (layer1_outputs(6836));
    layer2_outputs(6789) <= (layer1_outputs(9279)) xor (layer1_outputs(3117));
    layer2_outputs(6790) <= (layer1_outputs(2575)) or (layer1_outputs(5174));
    layer2_outputs(6791) <= not(layer1_outputs(4695));
    layer2_outputs(6792) <= not((layer1_outputs(7524)) and (layer1_outputs(5458)));
    layer2_outputs(6793) <= layer1_outputs(7287);
    layer2_outputs(6794) <= layer1_outputs(89);
    layer2_outputs(6795) <= layer1_outputs(2265);
    layer2_outputs(6796) <= not(layer1_outputs(4670));
    layer2_outputs(6797) <= layer1_outputs(6481);
    layer2_outputs(6798) <= not(layer1_outputs(388)) or (layer1_outputs(5770));
    layer2_outputs(6799) <= not(layer1_outputs(5619)) or (layer1_outputs(211));
    layer2_outputs(6800) <= layer1_outputs(2725);
    layer2_outputs(6801) <= (layer1_outputs(9801)) xor (layer1_outputs(3057));
    layer2_outputs(6802) <= (layer1_outputs(10)) and not (layer1_outputs(3650));
    layer2_outputs(6803) <= not(layer1_outputs(1966)) or (layer1_outputs(1781));
    layer2_outputs(6804) <= layer1_outputs(8705);
    layer2_outputs(6805) <= layer1_outputs(8515);
    layer2_outputs(6806) <= layer1_outputs(1979);
    layer2_outputs(6807) <= not(layer1_outputs(6365)) or (layer1_outputs(6338));
    layer2_outputs(6808) <= layer1_outputs(9847);
    layer2_outputs(6809) <= not(layer1_outputs(5895));
    layer2_outputs(6810) <= (layer1_outputs(2609)) and not (layer1_outputs(8899));
    layer2_outputs(6811) <= (layer1_outputs(1051)) or (layer1_outputs(7266));
    layer2_outputs(6812) <= layer1_outputs(10169);
    layer2_outputs(6813) <= (layer1_outputs(8580)) and not (layer1_outputs(5637));
    layer2_outputs(6814) <= not(layer1_outputs(4544)) or (layer1_outputs(9436));
    layer2_outputs(6815) <= layer1_outputs(2745);
    layer2_outputs(6816) <= layer1_outputs(107);
    layer2_outputs(6817) <= layer1_outputs(2978);
    layer2_outputs(6818) <= not(layer1_outputs(9355));
    layer2_outputs(6819) <= not(layer1_outputs(1231));
    layer2_outputs(6820) <= (layer1_outputs(8752)) xor (layer1_outputs(5561));
    layer2_outputs(6821) <= not(layer1_outputs(9153));
    layer2_outputs(6822) <= not(layer1_outputs(40));
    layer2_outputs(6823) <= not((layer1_outputs(5399)) or (layer1_outputs(1147)));
    layer2_outputs(6824) <= layer1_outputs(1830);
    layer2_outputs(6825) <= not((layer1_outputs(9187)) or (layer1_outputs(2807)));
    layer2_outputs(6826) <= '0';
    layer2_outputs(6827) <= layer1_outputs(9346);
    layer2_outputs(6828) <= not(layer1_outputs(2304));
    layer2_outputs(6829) <= not(layer1_outputs(6572));
    layer2_outputs(6830) <= not(layer1_outputs(8965));
    layer2_outputs(6831) <= layer1_outputs(67);
    layer2_outputs(6832) <= not(layer1_outputs(6251)) or (layer1_outputs(3032));
    layer2_outputs(6833) <= not(layer1_outputs(220)) or (layer1_outputs(2145));
    layer2_outputs(6834) <= not(layer1_outputs(6745));
    layer2_outputs(6835) <= (layer1_outputs(5722)) and not (layer1_outputs(6872));
    layer2_outputs(6836) <= layer1_outputs(1889);
    layer2_outputs(6837) <= not(layer1_outputs(1337)) or (layer1_outputs(10235));
    layer2_outputs(6838) <= layer1_outputs(3555);
    layer2_outputs(6839) <= (layer1_outputs(4442)) and not (layer1_outputs(6818));
    layer2_outputs(6840) <= not((layer1_outputs(4403)) or (layer1_outputs(6888)));
    layer2_outputs(6841) <= not((layer1_outputs(7604)) xor (layer1_outputs(8755)));
    layer2_outputs(6842) <= not(layer1_outputs(4883));
    layer2_outputs(6843) <= layer1_outputs(5133);
    layer2_outputs(6844) <= layer1_outputs(5699);
    layer2_outputs(6845) <= not(layer1_outputs(4797));
    layer2_outputs(6846) <= not((layer1_outputs(8025)) xor (layer1_outputs(1490)));
    layer2_outputs(6847) <= layer1_outputs(9203);
    layer2_outputs(6848) <= layer1_outputs(8204);
    layer2_outputs(6849) <= layer1_outputs(7279);
    layer2_outputs(6850) <= layer1_outputs(542);
    layer2_outputs(6851) <= layer1_outputs(3848);
    layer2_outputs(6852) <= (layer1_outputs(9008)) and not (layer1_outputs(1566));
    layer2_outputs(6853) <= not(layer1_outputs(4929));
    layer2_outputs(6854) <= layer1_outputs(3519);
    layer2_outputs(6855) <= not(layer1_outputs(6261));
    layer2_outputs(6856) <= (layer1_outputs(7228)) or (layer1_outputs(34));
    layer2_outputs(6857) <= layer1_outputs(6645);
    layer2_outputs(6858) <= not((layer1_outputs(5337)) or (layer1_outputs(714)));
    layer2_outputs(6859) <= not((layer1_outputs(3090)) xor (layer1_outputs(6521)));
    layer2_outputs(6860) <= not((layer1_outputs(322)) xor (layer1_outputs(3901)));
    layer2_outputs(6861) <= not((layer1_outputs(9435)) and (layer1_outputs(1823)));
    layer2_outputs(6862) <= (layer1_outputs(967)) and not (layer1_outputs(1139));
    layer2_outputs(6863) <= not((layer1_outputs(2355)) xor (layer1_outputs(1486)));
    layer2_outputs(6864) <= (layer1_outputs(2421)) and not (layer1_outputs(2829));
    layer2_outputs(6865) <= layer1_outputs(2783);
    layer2_outputs(6866) <= not(layer1_outputs(523));
    layer2_outputs(6867) <= '0';
    layer2_outputs(6868) <= not(layer1_outputs(9502)) or (layer1_outputs(6427));
    layer2_outputs(6869) <= not(layer1_outputs(4804)) or (layer1_outputs(8479));
    layer2_outputs(6870) <= (layer1_outputs(7797)) or (layer1_outputs(9700));
    layer2_outputs(6871) <= not((layer1_outputs(8379)) and (layer1_outputs(5567)));
    layer2_outputs(6872) <= not(layer1_outputs(4385));
    layer2_outputs(6873) <= not((layer1_outputs(8202)) and (layer1_outputs(5315)));
    layer2_outputs(6874) <= layer1_outputs(9670);
    layer2_outputs(6875) <= layer1_outputs(3752);
    layer2_outputs(6876) <= layer1_outputs(7053);
    layer2_outputs(6877) <= not((layer1_outputs(2235)) and (layer1_outputs(116)));
    layer2_outputs(6878) <= (layer1_outputs(9416)) and (layer1_outputs(6799));
    layer2_outputs(6879) <= not((layer1_outputs(4817)) xor (layer1_outputs(10018)));
    layer2_outputs(6880) <= not(layer1_outputs(2458)) or (layer1_outputs(3728));
    layer2_outputs(6881) <= (layer1_outputs(584)) and (layer1_outputs(6746));
    layer2_outputs(6882) <= (layer1_outputs(3817)) and (layer1_outputs(2280));
    layer2_outputs(6883) <= not((layer1_outputs(6679)) xor (layer1_outputs(9163)));
    layer2_outputs(6884) <= (layer1_outputs(3445)) or (layer1_outputs(7771));
    layer2_outputs(6885) <= (layer1_outputs(8397)) or (layer1_outputs(469));
    layer2_outputs(6886) <= (layer1_outputs(1264)) and not (layer1_outputs(2038));
    layer2_outputs(6887) <= (layer1_outputs(6482)) xor (layer1_outputs(1567));
    layer2_outputs(6888) <= layer1_outputs(5516);
    layer2_outputs(6889) <= (layer1_outputs(9766)) and not (layer1_outputs(7198));
    layer2_outputs(6890) <= layer1_outputs(2106);
    layer2_outputs(6891) <= layer1_outputs(965);
    layer2_outputs(6892) <= (layer1_outputs(2891)) and (layer1_outputs(3553));
    layer2_outputs(6893) <= not(layer1_outputs(2032));
    layer2_outputs(6894) <= layer1_outputs(5127);
    layer2_outputs(6895) <= not(layer1_outputs(1005));
    layer2_outputs(6896) <= (layer1_outputs(10073)) and not (layer1_outputs(5659));
    layer2_outputs(6897) <= not(layer1_outputs(7472));
    layer2_outputs(6898) <= (layer1_outputs(8988)) or (layer1_outputs(6771));
    layer2_outputs(6899) <= (layer1_outputs(4782)) xor (layer1_outputs(4989));
    layer2_outputs(6900) <= not((layer1_outputs(6394)) xor (layer1_outputs(1544)));
    layer2_outputs(6901) <= not(layer1_outputs(922)) or (layer1_outputs(7672));
    layer2_outputs(6902) <= not(layer1_outputs(2209)) or (layer1_outputs(6079));
    layer2_outputs(6903) <= layer1_outputs(1440);
    layer2_outputs(6904) <= (layer1_outputs(5212)) and not (layer1_outputs(3898));
    layer2_outputs(6905) <= (layer1_outputs(6163)) and not (layer1_outputs(9825));
    layer2_outputs(6906) <= (layer1_outputs(2564)) and (layer1_outputs(1235));
    layer2_outputs(6907) <= not(layer1_outputs(7141));
    layer2_outputs(6908) <= not(layer1_outputs(4115)) or (layer1_outputs(2042));
    layer2_outputs(6909) <= not(layer1_outputs(8096));
    layer2_outputs(6910) <= not(layer1_outputs(5095));
    layer2_outputs(6911) <= not(layer1_outputs(1534));
    layer2_outputs(6912) <= (layer1_outputs(5012)) xor (layer1_outputs(6719));
    layer2_outputs(6913) <= layer1_outputs(6274);
    layer2_outputs(6914) <= not(layer1_outputs(5677));
    layer2_outputs(6915) <= (layer1_outputs(7600)) or (layer1_outputs(9712));
    layer2_outputs(6916) <= layer1_outputs(3347);
    layer2_outputs(6917) <= (layer1_outputs(9445)) and (layer1_outputs(5053));
    layer2_outputs(6918) <= layer1_outputs(3536);
    layer2_outputs(6919) <= not(layer1_outputs(470)) or (layer1_outputs(8824));
    layer2_outputs(6920) <= not((layer1_outputs(82)) xor (layer1_outputs(6430)));
    layer2_outputs(6921) <= not((layer1_outputs(3757)) and (layer1_outputs(1332)));
    layer2_outputs(6922) <= (layer1_outputs(3980)) and not (layer1_outputs(5607));
    layer2_outputs(6923) <= layer1_outputs(6728);
    layer2_outputs(6924) <= not(layer1_outputs(1512));
    layer2_outputs(6925) <= layer1_outputs(7975);
    layer2_outputs(6926) <= '0';
    layer2_outputs(6927) <= (layer1_outputs(7839)) xor (layer1_outputs(7246));
    layer2_outputs(6928) <= not(layer1_outputs(1020));
    layer2_outputs(6929) <= (layer1_outputs(4382)) xor (layer1_outputs(9060));
    layer2_outputs(6930) <= not((layer1_outputs(4566)) and (layer1_outputs(6375)));
    layer2_outputs(6931) <= layer1_outputs(8212);
    layer2_outputs(6932) <= (layer1_outputs(6433)) and not (layer1_outputs(9357));
    layer2_outputs(6933) <= not((layer1_outputs(7150)) xor (layer1_outputs(5772)));
    layer2_outputs(6934) <= (layer1_outputs(5786)) and not (layer1_outputs(108));
    layer2_outputs(6935) <= not((layer1_outputs(16)) or (layer1_outputs(6032)));
    layer2_outputs(6936) <= not(layer1_outputs(4048));
    layer2_outputs(6937) <= (layer1_outputs(6725)) and not (layer1_outputs(5488));
    layer2_outputs(6938) <= not(layer1_outputs(4364));
    layer2_outputs(6939) <= (layer1_outputs(818)) xor (layer1_outputs(2914));
    layer2_outputs(6940) <= not(layer1_outputs(2098));
    layer2_outputs(6941) <= not(layer1_outputs(9546));
    layer2_outputs(6942) <= not((layer1_outputs(3277)) or (layer1_outputs(6119)));
    layer2_outputs(6943) <= not(layer1_outputs(4152)) or (layer1_outputs(853));
    layer2_outputs(6944) <= '1';
    layer2_outputs(6945) <= not((layer1_outputs(9097)) or (layer1_outputs(2791)));
    layer2_outputs(6946) <= not(layer1_outputs(9367));
    layer2_outputs(6947) <= not(layer1_outputs(8337));
    layer2_outputs(6948) <= '1';
    layer2_outputs(6949) <= not((layer1_outputs(6115)) and (layer1_outputs(5106)));
    layer2_outputs(6950) <= layer1_outputs(8452);
    layer2_outputs(6951) <= (layer1_outputs(8140)) xor (layer1_outputs(1069));
    layer2_outputs(6952) <= not(layer1_outputs(8297)) or (layer1_outputs(1385));
    layer2_outputs(6953) <= not(layer1_outputs(3739));
    layer2_outputs(6954) <= not((layer1_outputs(2593)) or (layer1_outputs(3951)));
    layer2_outputs(6955) <= not(layer1_outputs(572));
    layer2_outputs(6956) <= (layer1_outputs(9458)) and not (layer1_outputs(354));
    layer2_outputs(6957) <= (layer1_outputs(8645)) xor (layer1_outputs(3929));
    layer2_outputs(6958) <= '1';
    layer2_outputs(6959) <= (layer1_outputs(8364)) xor (layer1_outputs(8148));
    layer2_outputs(6960) <= layer1_outputs(4080);
    layer2_outputs(6961) <= not(layer1_outputs(7663));
    layer2_outputs(6962) <= not(layer1_outputs(9444)) or (layer1_outputs(7998));
    layer2_outputs(6963) <= layer1_outputs(4580);
    layer2_outputs(6964) <= (layer1_outputs(4928)) xor (layer1_outputs(6716));
    layer2_outputs(6965) <= not(layer1_outputs(72)) or (layer1_outputs(4363));
    layer2_outputs(6966) <= not((layer1_outputs(5730)) or (layer1_outputs(7086)));
    layer2_outputs(6967) <= not(layer1_outputs(6607)) or (layer1_outputs(5436));
    layer2_outputs(6968) <= (layer1_outputs(3190)) and (layer1_outputs(4470));
    layer2_outputs(6969) <= not(layer1_outputs(2799));
    layer2_outputs(6970) <= layer1_outputs(3809);
    layer2_outputs(6971) <= not((layer1_outputs(6897)) and (layer1_outputs(6333)));
    layer2_outputs(6972) <= not(layer1_outputs(5967));
    layer2_outputs(6973) <= (layer1_outputs(78)) and not (layer1_outputs(3845));
    layer2_outputs(6974) <= layer1_outputs(7916);
    layer2_outputs(6975) <= not(layer1_outputs(8924)) or (layer1_outputs(1162));
    layer2_outputs(6976) <= not(layer1_outputs(3082)) or (layer1_outputs(6201));
    layer2_outputs(6977) <= (layer1_outputs(2287)) xor (layer1_outputs(9139));
    layer2_outputs(6978) <= not(layer1_outputs(1599));
    layer2_outputs(6979) <= (layer1_outputs(184)) or (layer1_outputs(5690));
    layer2_outputs(6980) <= not(layer1_outputs(769));
    layer2_outputs(6981) <= not(layer1_outputs(6365));
    layer2_outputs(6982) <= layer1_outputs(10165);
    layer2_outputs(6983) <= (layer1_outputs(4833)) xor (layer1_outputs(9340));
    layer2_outputs(6984) <= layer1_outputs(6087);
    layer2_outputs(6985) <= not(layer1_outputs(1151)) or (layer1_outputs(2607));
    layer2_outputs(6986) <= not((layer1_outputs(8111)) and (layer1_outputs(3376)));
    layer2_outputs(6987) <= not((layer1_outputs(8523)) and (layer1_outputs(5195)));
    layer2_outputs(6988) <= not(layer1_outputs(9606));
    layer2_outputs(6989) <= not((layer1_outputs(1085)) xor (layer1_outputs(3724)));
    layer2_outputs(6990) <= layer1_outputs(5485);
    layer2_outputs(6991) <= (layer1_outputs(4650)) and (layer1_outputs(8644));
    layer2_outputs(6992) <= not(layer1_outputs(3586));
    layer2_outputs(6993) <= not(layer1_outputs(7055));
    layer2_outputs(6994) <= (layer1_outputs(1485)) and not (layer1_outputs(3616));
    layer2_outputs(6995) <= not(layer1_outputs(3219));
    layer2_outputs(6996) <= layer1_outputs(839);
    layer2_outputs(6997) <= not(layer1_outputs(7440)) or (layer1_outputs(4613));
    layer2_outputs(6998) <= (layer1_outputs(1643)) or (layer1_outputs(428));
    layer2_outputs(6999) <= not((layer1_outputs(4861)) and (layer1_outputs(920)));
    layer2_outputs(7000) <= (layer1_outputs(4395)) and not (layer1_outputs(2462));
    layer2_outputs(7001) <= not(layer1_outputs(9844));
    layer2_outputs(7002) <= not(layer1_outputs(5240));
    layer2_outputs(7003) <= (layer1_outputs(3173)) or (layer1_outputs(5119));
    layer2_outputs(7004) <= not((layer1_outputs(2642)) xor (layer1_outputs(9251)));
    layer2_outputs(7005) <= not(layer1_outputs(5545));
    layer2_outputs(7006) <= not(layer1_outputs(5834));
    layer2_outputs(7007) <= layer1_outputs(226);
    layer2_outputs(7008) <= (layer1_outputs(5306)) and not (layer1_outputs(7506));
    layer2_outputs(7009) <= not(layer1_outputs(8788)) or (layer1_outputs(3624));
    layer2_outputs(7010) <= layer1_outputs(3995);
    layer2_outputs(7011) <= (layer1_outputs(9781)) xor (layer1_outputs(6540));
    layer2_outputs(7012) <= not(layer1_outputs(547));
    layer2_outputs(7013) <= (layer1_outputs(3627)) and not (layer1_outputs(8460));
    layer2_outputs(7014) <= not((layer1_outputs(2489)) xor (layer1_outputs(1783)));
    layer2_outputs(7015) <= not((layer1_outputs(4810)) xor (layer1_outputs(9375)));
    layer2_outputs(7016) <= not(layer1_outputs(2506)) or (layer1_outputs(9958));
    layer2_outputs(7017) <= (layer1_outputs(5217)) and not (layer1_outputs(4653));
    layer2_outputs(7018) <= layer1_outputs(8340);
    layer2_outputs(7019) <= layer1_outputs(8214);
    layer2_outputs(7020) <= (layer1_outputs(4735)) and (layer1_outputs(2329));
    layer2_outputs(7021) <= not(layer1_outputs(2559));
    layer2_outputs(7022) <= not(layer1_outputs(10210));
    layer2_outputs(7023) <= not(layer1_outputs(4438)) or (layer1_outputs(2800));
    layer2_outputs(7024) <= layer1_outputs(7648);
    layer2_outputs(7025) <= not((layer1_outputs(5269)) or (layer1_outputs(258)));
    layer2_outputs(7026) <= not(layer1_outputs(8232));
    layer2_outputs(7027) <= (layer1_outputs(3082)) and not (layer1_outputs(3839));
    layer2_outputs(7028) <= layer1_outputs(7067);
    layer2_outputs(7029) <= not(layer1_outputs(9169));
    layer2_outputs(7030) <= not((layer1_outputs(3768)) xor (layer1_outputs(4493)));
    layer2_outputs(7031) <= not(layer1_outputs(9526)) or (layer1_outputs(5596));
    layer2_outputs(7032) <= (layer1_outputs(3993)) or (layer1_outputs(5527));
    layer2_outputs(7033) <= not((layer1_outputs(8467)) and (layer1_outputs(3592)));
    layer2_outputs(7034) <= not(layer1_outputs(4646));
    layer2_outputs(7035) <= not(layer1_outputs(3994));
    layer2_outputs(7036) <= not(layer1_outputs(7490));
    layer2_outputs(7037) <= (layer1_outputs(4145)) and not (layer1_outputs(1443));
    layer2_outputs(7038) <= not(layer1_outputs(6256));
    layer2_outputs(7039) <= layer1_outputs(3868);
    layer2_outputs(7040) <= layer1_outputs(8783);
    layer2_outputs(7041) <= layer1_outputs(4085);
    layer2_outputs(7042) <= not(layer1_outputs(1850)) or (layer1_outputs(2180));
    layer2_outputs(7043) <= not(layer1_outputs(1268));
    layer2_outputs(7044) <= not((layer1_outputs(6325)) xor (layer1_outputs(7025)));
    layer2_outputs(7045) <= not((layer1_outputs(7895)) xor (layer1_outputs(1024)));
    layer2_outputs(7046) <= not((layer1_outputs(6307)) xor (layer1_outputs(3656)));
    layer2_outputs(7047) <= not(layer1_outputs(6428));
    layer2_outputs(7048) <= not(layer1_outputs(3852));
    layer2_outputs(7049) <= not(layer1_outputs(1260));
    layer2_outputs(7050) <= not(layer1_outputs(3841));
    layer2_outputs(7051) <= layer1_outputs(1200);
    layer2_outputs(7052) <= layer1_outputs(323);
    layer2_outputs(7053) <= not((layer1_outputs(2011)) or (layer1_outputs(1358)));
    layer2_outputs(7054) <= not((layer1_outputs(8480)) and (layer1_outputs(1363)));
    layer2_outputs(7055) <= not((layer1_outputs(8834)) xor (layer1_outputs(6933)));
    layer2_outputs(7056) <= not(layer1_outputs(3510)) or (layer1_outputs(1852));
    layer2_outputs(7057) <= layer1_outputs(7051);
    layer2_outputs(7058) <= not((layer1_outputs(6414)) xor (layer1_outputs(1321)));
    layer2_outputs(7059) <= (layer1_outputs(8146)) and not (layer1_outputs(730));
    layer2_outputs(7060) <= not(layer1_outputs(6828));
    layer2_outputs(7061) <= (layer1_outputs(10100)) and not (layer1_outputs(5186));
    layer2_outputs(7062) <= not(layer1_outputs(1986));
    layer2_outputs(7063) <= (layer1_outputs(9485)) and not (layer1_outputs(3707));
    layer2_outputs(7064) <= (layer1_outputs(4425)) and not (layer1_outputs(5877));
    layer2_outputs(7065) <= not(layer1_outputs(10162));
    layer2_outputs(7066) <= layer1_outputs(944);
    layer2_outputs(7067) <= not((layer1_outputs(1910)) and (layer1_outputs(7753)));
    layer2_outputs(7068) <= layer1_outputs(4535);
    layer2_outputs(7069) <= not(layer1_outputs(8833));
    layer2_outputs(7070) <= not(layer1_outputs(5777)) or (layer1_outputs(4689));
    layer2_outputs(7071) <= not(layer1_outputs(1091));
    layer2_outputs(7072) <= not((layer1_outputs(9552)) or (layer1_outputs(45)));
    layer2_outputs(7073) <= (layer1_outputs(6086)) xor (layer1_outputs(819));
    layer2_outputs(7074) <= not(layer1_outputs(23));
    layer2_outputs(7075) <= (layer1_outputs(4464)) and not (layer1_outputs(9909));
    layer2_outputs(7076) <= (layer1_outputs(1519)) xor (layer1_outputs(5375));
    layer2_outputs(7077) <= layer1_outputs(2135);
    layer2_outputs(7078) <= not(layer1_outputs(1211));
    layer2_outputs(7079) <= (layer1_outputs(8629)) and not (layer1_outputs(5439));
    layer2_outputs(7080) <= layer1_outputs(4024);
    layer2_outputs(7081) <= not(layer1_outputs(7318));
    layer2_outputs(7082) <= not(layer1_outputs(4270));
    layer2_outputs(7083) <= not((layer1_outputs(188)) or (layer1_outputs(7653)));
    layer2_outputs(7084) <= not(layer1_outputs(3488)) or (layer1_outputs(5678));
    layer2_outputs(7085) <= not(layer1_outputs(4737)) or (layer1_outputs(3018));
    layer2_outputs(7086) <= (layer1_outputs(1868)) xor (layer1_outputs(6216));
    layer2_outputs(7087) <= not(layer1_outputs(8244));
    layer2_outputs(7088) <= layer1_outputs(1831);
    layer2_outputs(7089) <= (layer1_outputs(7647)) and not (layer1_outputs(5674));
    layer2_outputs(7090) <= layer1_outputs(8795);
    layer2_outputs(7091) <= not(layer1_outputs(4507));
    layer2_outputs(7092) <= not(layer1_outputs(6575)) or (layer1_outputs(6539));
    layer2_outputs(7093) <= layer1_outputs(7525);
    layer2_outputs(7094) <= (layer1_outputs(8623)) or (layer1_outputs(5840));
    layer2_outputs(7095) <= (layer1_outputs(4844)) and not (layer1_outputs(7421));
    layer2_outputs(7096) <= layer1_outputs(8632);
    layer2_outputs(7097) <= not((layer1_outputs(911)) and (layer1_outputs(2901)));
    layer2_outputs(7098) <= (layer1_outputs(3116)) xor (layer1_outputs(3312));
    layer2_outputs(7099) <= layer1_outputs(556);
    layer2_outputs(7100) <= not(layer1_outputs(6470)) or (layer1_outputs(9839));
    layer2_outputs(7101) <= not((layer1_outputs(5221)) or (layer1_outputs(1158)));
    layer2_outputs(7102) <= not(layer1_outputs(10231)) or (layer1_outputs(7215));
    layer2_outputs(7103) <= not(layer1_outputs(4072));
    layer2_outputs(7104) <= not((layer1_outputs(4003)) and (layer1_outputs(4561)));
    layer2_outputs(7105) <= (layer1_outputs(1991)) or (layer1_outputs(5099));
    layer2_outputs(7106) <= layer1_outputs(9486);
    layer2_outputs(7107) <= not(layer1_outputs(7312)) or (layer1_outputs(4569));
    layer2_outputs(7108) <= not(layer1_outputs(8677)) or (layer1_outputs(9961));
    layer2_outputs(7109) <= (layer1_outputs(9354)) xor (layer1_outputs(5191));
    layer2_outputs(7110) <= layer1_outputs(8882);
    layer2_outputs(7111) <= layer1_outputs(5438);
    layer2_outputs(7112) <= not((layer1_outputs(896)) and (layer1_outputs(7569)));
    layer2_outputs(7113) <= layer1_outputs(10160);
    layer2_outputs(7114) <= not(layer1_outputs(697));
    layer2_outputs(7115) <= not((layer1_outputs(9974)) xor (layer1_outputs(5287)));
    layer2_outputs(7116) <= not(layer1_outputs(4743));
    layer2_outputs(7117) <= (layer1_outputs(6009)) and (layer1_outputs(9248));
    layer2_outputs(7118) <= not(layer1_outputs(7764)) or (layer1_outputs(8741));
    layer2_outputs(7119) <= (layer1_outputs(3475)) and not (layer1_outputs(3304));
    layer2_outputs(7120) <= not(layer1_outputs(3467));
    layer2_outputs(7121) <= layer1_outputs(1837);
    layer2_outputs(7122) <= not(layer1_outputs(3886));
    layer2_outputs(7123) <= (layer1_outputs(5377)) or (layer1_outputs(4130));
    layer2_outputs(7124) <= not(layer1_outputs(1639));
    layer2_outputs(7125) <= layer1_outputs(1805);
    layer2_outputs(7126) <= '0';
    layer2_outputs(7127) <= not(layer1_outputs(8476));
    layer2_outputs(7128) <= layer1_outputs(7212);
    layer2_outputs(7129) <= (layer1_outputs(4428)) and not (layer1_outputs(3787));
    layer2_outputs(7130) <= (layer1_outputs(9195)) and not (layer1_outputs(7884));
    layer2_outputs(7131) <= not((layer1_outputs(5553)) and (layer1_outputs(2931)));
    layer2_outputs(7132) <= layer1_outputs(1594);
    layer2_outputs(7133) <= layer1_outputs(7859);
    layer2_outputs(7134) <= layer1_outputs(564);
    layer2_outputs(7135) <= layer1_outputs(9805);
    layer2_outputs(7136) <= not(layer1_outputs(4368));
    layer2_outputs(7137) <= not(layer1_outputs(4421));
    layer2_outputs(7138) <= layer1_outputs(6254);
    layer2_outputs(7139) <= not(layer1_outputs(1980)) or (layer1_outputs(1150));
    layer2_outputs(7140) <= not(layer1_outputs(2341));
    layer2_outputs(7141) <= not(layer1_outputs(1091));
    layer2_outputs(7142) <= not((layer1_outputs(7567)) or (layer1_outputs(5523)));
    layer2_outputs(7143) <= layer1_outputs(6801);
    layer2_outputs(7144) <= (layer1_outputs(5341)) and not (layer1_outputs(1464));
    layer2_outputs(7145) <= not(layer1_outputs(8923));
    layer2_outputs(7146) <= (layer1_outputs(1248)) and not (layer1_outputs(7692));
    layer2_outputs(7147) <= (layer1_outputs(7141)) xor (layer1_outputs(4986));
    layer2_outputs(7148) <= (layer1_outputs(6060)) and not (layer1_outputs(6710));
    layer2_outputs(7149) <= not(layer1_outputs(1361));
    layer2_outputs(7150) <= layer1_outputs(1127);
    layer2_outputs(7151) <= (layer1_outputs(1222)) and not (layer1_outputs(1028));
    layer2_outputs(7152) <= not((layer1_outputs(1238)) xor (layer1_outputs(5456)));
    layer2_outputs(7153) <= layer1_outputs(7397);
    layer2_outputs(7154) <= layer1_outputs(9376);
    layer2_outputs(7155) <= not((layer1_outputs(408)) or (layer1_outputs(9421)));
    layer2_outputs(7156) <= (layer1_outputs(9937)) or (layer1_outputs(3970));
    layer2_outputs(7157) <= not((layer1_outputs(7845)) xor (layer1_outputs(7326)));
    layer2_outputs(7158) <= not(layer1_outputs(2371)) or (layer1_outputs(7444));
    layer2_outputs(7159) <= (layer1_outputs(5447)) xor (layer1_outputs(7192));
    layer2_outputs(7160) <= not(layer1_outputs(8065));
    layer2_outputs(7161) <= not(layer1_outputs(1148));
    layer2_outputs(7162) <= not(layer1_outputs(3403));
    layer2_outputs(7163) <= not((layer1_outputs(4286)) and (layer1_outputs(7782)));
    layer2_outputs(7164) <= (layer1_outputs(4765)) xor (layer1_outputs(3149));
    layer2_outputs(7165) <= not(layer1_outputs(4398)) or (layer1_outputs(1107));
    layer2_outputs(7166) <= not(layer1_outputs(7750));
    layer2_outputs(7167) <= not(layer1_outputs(6804));
    layer2_outputs(7168) <= not((layer1_outputs(2173)) or (layer1_outputs(5478)));
    layer2_outputs(7169) <= not(layer1_outputs(7348));
    layer2_outputs(7170) <= '1';
    layer2_outputs(7171) <= '1';
    layer2_outputs(7172) <= not(layer1_outputs(4912)) or (layer1_outputs(9754));
    layer2_outputs(7173) <= not(layer1_outputs(4502));
    layer2_outputs(7174) <= not(layer1_outputs(1731));
    layer2_outputs(7175) <= (layer1_outputs(6318)) and not (layer1_outputs(4543));
    layer2_outputs(7176) <= not(layer1_outputs(4554)) or (layer1_outputs(5018));
    layer2_outputs(7177) <= not(layer1_outputs(1522));
    layer2_outputs(7178) <= (layer1_outputs(1138)) and not (layer1_outputs(2479));
    layer2_outputs(7179) <= not(layer1_outputs(9453)) or (layer1_outputs(703));
    layer2_outputs(7180) <= layer1_outputs(6180);
    layer2_outputs(7181) <= layer1_outputs(6014);
    layer2_outputs(7182) <= not((layer1_outputs(4193)) xor (layer1_outputs(7295)));
    layer2_outputs(7183) <= layer1_outputs(1124);
    layer2_outputs(7184) <= (layer1_outputs(4379)) xor (layer1_outputs(372));
    layer2_outputs(7185) <= '0';
    layer2_outputs(7186) <= not((layer1_outputs(8433)) and (layer1_outputs(4943)));
    layer2_outputs(7187) <= not(layer1_outputs(4293));
    layer2_outputs(7188) <= layer1_outputs(5353);
    layer2_outputs(7189) <= '1';
    layer2_outputs(7190) <= (layer1_outputs(4889)) and not (layer1_outputs(3216));
    layer2_outputs(7191) <= (layer1_outputs(8420)) and not (layer1_outputs(4376));
    layer2_outputs(7192) <= layer1_outputs(1367);
    layer2_outputs(7193) <= not(layer1_outputs(165));
    layer2_outputs(7194) <= (layer1_outputs(9258)) and not (layer1_outputs(936));
    layer2_outputs(7195) <= (layer1_outputs(1376)) and not (layer1_outputs(8984));
    layer2_outputs(7196) <= (layer1_outputs(259)) xor (layer1_outputs(216));
    layer2_outputs(7197) <= (layer1_outputs(7571)) and not (layer1_outputs(1307));
    layer2_outputs(7198) <= layer1_outputs(9744);
    layer2_outputs(7199) <= layer1_outputs(5386);
    layer2_outputs(7200) <= layer1_outputs(849);
    layer2_outputs(7201) <= layer1_outputs(4511);
    layer2_outputs(7202) <= layer1_outputs(2506);
    layer2_outputs(7203) <= (layer1_outputs(3516)) and not (layer1_outputs(2507));
    layer2_outputs(7204) <= not(layer1_outputs(8868)) or (layer1_outputs(9309));
    layer2_outputs(7205) <= (layer1_outputs(405)) and not (layer1_outputs(8674));
    layer2_outputs(7206) <= not((layer1_outputs(1563)) xor (layer1_outputs(6197)));
    layer2_outputs(7207) <= not(layer1_outputs(6359));
    layer2_outputs(7208) <= '1';
    layer2_outputs(7209) <= layer1_outputs(134);
    layer2_outputs(7210) <= (layer1_outputs(7410)) or (layer1_outputs(136));
    layer2_outputs(7211) <= not(layer1_outputs(2927));
    layer2_outputs(7212) <= not(layer1_outputs(9833));
    layer2_outputs(7213) <= layer1_outputs(5950);
    layer2_outputs(7214) <= not(layer1_outputs(2898));
    layer2_outputs(7215) <= not(layer1_outputs(195));
    layer2_outputs(7216) <= (layer1_outputs(3295)) and not (layer1_outputs(396));
    layer2_outputs(7217) <= layer1_outputs(2447);
    layer2_outputs(7218) <= (layer1_outputs(3612)) and not (layer1_outputs(9345));
    layer2_outputs(7219) <= layer1_outputs(4312);
    layer2_outputs(7220) <= not(layer1_outputs(5636));
    layer2_outputs(7221) <= not(layer1_outputs(1005));
    layer2_outputs(7222) <= layer1_outputs(3079);
    layer2_outputs(7223) <= not(layer1_outputs(9344));
    layer2_outputs(7224) <= not(layer1_outputs(10221)) or (layer1_outputs(6949));
    layer2_outputs(7225) <= not(layer1_outputs(1595));
    layer2_outputs(7226) <= '1';
    layer2_outputs(7227) <= layer1_outputs(9240);
    layer2_outputs(7228) <= layer1_outputs(2278);
    layer2_outputs(7229) <= '1';
    layer2_outputs(7230) <= not((layer1_outputs(8285)) or (layer1_outputs(9668)));
    layer2_outputs(7231) <= not(layer1_outputs(5002));
    layer2_outputs(7232) <= not((layer1_outputs(1126)) xor (layer1_outputs(5208)));
    layer2_outputs(7233) <= layer1_outputs(109);
    layer2_outputs(7234) <= not((layer1_outputs(1539)) xor (layer1_outputs(1639)));
    layer2_outputs(7235) <= not((layer1_outputs(1558)) xor (layer1_outputs(9462)));
    layer2_outputs(7236) <= (layer1_outputs(8497)) xor (layer1_outputs(1307));
    layer2_outputs(7237) <= (layer1_outputs(1829)) and (layer1_outputs(8079));
    layer2_outputs(7238) <= (layer1_outputs(2869)) or (layer1_outputs(9391));
    layer2_outputs(7239) <= not((layer1_outputs(2639)) xor (layer1_outputs(3434)));
    layer2_outputs(7240) <= (layer1_outputs(6400)) and (layer1_outputs(9530));
    layer2_outputs(7241) <= (layer1_outputs(5500)) and (layer1_outputs(5733));
    layer2_outputs(7242) <= not((layer1_outputs(5277)) xor (layer1_outputs(7608)));
    layer2_outputs(7243) <= layer1_outputs(3913);
    layer2_outputs(7244) <= layer1_outputs(3433);
    layer2_outputs(7245) <= (layer1_outputs(2335)) and not (layer1_outputs(3168));
    layer2_outputs(7246) <= not((layer1_outputs(8188)) and (layer1_outputs(6780)));
    layer2_outputs(7247) <= not((layer1_outputs(3074)) or (layer1_outputs(163)));
    layer2_outputs(7248) <= layer1_outputs(2439);
    layer2_outputs(7249) <= not(layer1_outputs(8728));
    layer2_outputs(7250) <= (layer1_outputs(4327)) xor (layer1_outputs(899));
    layer2_outputs(7251) <= layer1_outputs(2025);
    layer2_outputs(7252) <= (layer1_outputs(1312)) xor (layer1_outputs(3803));
    layer2_outputs(7253) <= layer1_outputs(5114);
    layer2_outputs(7254) <= not((layer1_outputs(1294)) xor (layer1_outputs(2693)));
    layer2_outputs(7255) <= not(layer1_outputs(6601));
    layer2_outputs(7256) <= layer1_outputs(9154);
    layer2_outputs(7257) <= (layer1_outputs(6648)) and not (layer1_outputs(9303));
    layer2_outputs(7258) <= layer1_outputs(4386);
    layer2_outputs(7259) <= not(layer1_outputs(831)) or (layer1_outputs(4504));
    layer2_outputs(7260) <= (layer1_outputs(8282)) and not (layer1_outputs(3802));
    layer2_outputs(7261) <= (layer1_outputs(1726)) and not (layer1_outputs(3746));
    layer2_outputs(7262) <= (layer1_outputs(4641)) and (layer1_outputs(4936));
    layer2_outputs(7263) <= (layer1_outputs(8862)) and not (layer1_outputs(781));
    layer2_outputs(7264) <= layer1_outputs(3457);
    layer2_outputs(7265) <= (layer1_outputs(4003)) and not (layer1_outputs(8892));
    layer2_outputs(7266) <= not(layer1_outputs(9155));
    layer2_outputs(7267) <= not(layer1_outputs(7386));
    layer2_outputs(7268) <= layer1_outputs(8221);
    layer2_outputs(7269) <= layer1_outputs(7776);
    layer2_outputs(7270) <= not((layer1_outputs(3499)) xor (layer1_outputs(2916)));
    layer2_outputs(7271) <= (layer1_outputs(9490)) and not (layer1_outputs(8628));
    layer2_outputs(7272) <= layer1_outputs(4443);
    layer2_outputs(7273) <= not((layer1_outputs(180)) or (layer1_outputs(6568)));
    layer2_outputs(7274) <= not((layer1_outputs(7550)) xor (layer1_outputs(4335)));
    layer2_outputs(7275) <= not(layer1_outputs(4088));
    layer2_outputs(7276) <= (layer1_outputs(8281)) and (layer1_outputs(3491));
    layer2_outputs(7277) <= not(layer1_outputs(8435));
    layer2_outputs(7278) <= not(layer1_outputs(3221)) or (layer1_outputs(2242));
    layer2_outputs(7279) <= (layer1_outputs(6533)) and not (layer1_outputs(10225));
    layer2_outputs(7280) <= (layer1_outputs(4039)) xor (layer1_outputs(7250));
    layer2_outputs(7281) <= not((layer1_outputs(6122)) or (layer1_outputs(10233)));
    layer2_outputs(7282) <= not(layer1_outputs(1365)) or (layer1_outputs(2013));
    layer2_outputs(7283) <= (layer1_outputs(5129)) xor (layer1_outputs(5886));
    layer2_outputs(7284) <= layer1_outputs(2025);
    layer2_outputs(7285) <= (layer1_outputs(7179)) and not (layer1_outputs(9793));
    layer2_outputs(7286) <= not(layer1_outputs(2496)) or (layer1_outputs(8655));
    layer2_outputs(7287) <= not(layer1_outputs(5374));
    layer2_outputs(7288) <= layer1_outputs(4153);
    layer2_outputs(7289) <= not(layer1_outputs(5061)) or (layer1_outputs(1271));
    layer2_outputs(7290) <= (layer1_outputs(3601)) and (layer1_outputs(8978));
    layer2_outputs(7291) <= not(layer1_outputs(6978)) or (layer1_outputs(8457));
    layer2_outputs(7292) <= (layer1_outputs(1171)) and not (layer1_outputs(8408));
    layer2_outputs(7293) <= not((layer1_outputs(5844)) xor (layer1_outputs(98)));
    layer2_outputs(7294) <= not((layer1_outputs(493)) or (layer1_outputs(4760)));
    layer2_outputs(7295) <= not(layer1_outputs(2729));
    layer2_outputs(7296) <= not(layer1_outputs(8587)) or (layer1_outputs(1505));
    layer2_outputs(7297) <= layer1_outputs(4973);
    layer2_outputs(7298) <= layer1_outputs(7693);
    layer2_outputs(7299) <= not(layer1_outputs(1992));
    layer2_outputs(7300) <= not((layer1_outputs(9256)) and (layer1_outputs(145)));
    layer2_outputs(7301) <= not((layer1_outputs(5557)) and (layer1_outputs(3046)));
    layer2_outputs(7302) <= not(layer1_outputs(8770)) or (layer1_outputs(4956));
    layer2_outputs(7303) <= (layer1_outputs(7928)) and not (layer1_outputs(5480));
    layer2_outputs(7304) <= (layer1_outputs(6691)) and not (layer1_outputs(1647));
    layer2_outputs(7305) <= not((layer1_outputs(6673)) xor (layer1_outputs(7982)));
    layer2_outputs(7306) <= layer1_outputs(10089);
    layer2_outputs(7307) <= not(layer1_outputs(4704));
    layer2_outputs(7308) <= (layer1_outputs(9253)) and not (layer1_outputs(8631));
    layer2_outputs(7309) <= not(layer1_outputs(6786));
    layer2_outputs(7310) <= layer1_outputs(6060);
    layer2_outputs(7311) <= layer1_outputs(881);
    layer2_outputs(7312) <= layer1_outputs(8744);
    layer2_outputs(7313) <= layer1_outputs(1004);
    layer2_outputs(7314) <= (layer1_outputs(7985)) xor (layer1_outputs(7200));
    layer2_outputs(7315) <= not(layer1_outputs(5924));
    layer2_outputs(7316) <= not(layer1_outputs(9088));
    layer2_outputs(7317) <= not(layer1_outputs(2157));
    layer2_outputs(7318) <= not(layer1_outputs(1100));
    layer2_outputs(7319) <= not(layer1_outputs(7534));
    layer2_outputs(7320) <= layer1_outputs(9494);
    layer2_outputs(7321) <= layer1_outputs(1069);
    layer2_outputs(7322) <= not(layer1_outputs(4165));
    layer2_outputs(7323) <= (layer1_outputs(587)) and (layer1_outputs(2747));
    layer2_outputs(7324) <= not(layer1_outputs(3317));
    layer2_outputs(7325) <= layer1_outputs(6346);
    layer2_outputs(7326) <= not(layer1_outputs(1976));
    layer2_outputs(7327) <= not(layer1_outputs(7801));
    layer2_outputs(7328) <= not(layer1_outputs(6134));
    layer2_outputs(7329) <= layer1_outputs(2008);
    layer2_outputs(7330) <= (layer1_outputs(7823)) xor (layer1_outputs(5068));
    layer2_outputs(7331) <= (layer1_outputs(6640)) and not (layer1_outputs(5660));
    layer2_outputs(7332) <= (layer1_outputs(4579)) and not (layer1_outputs(2712));
    layer2_outputs(7333) <= not(layer1_outputs(4516)) or (layer1_outputs(7204));
    layer2_outputs(7334) <= layer1_outputs(1646);
    layer2_outputs(7335) <= not(layer1_outputs(7911));
    layer2_outputs(7336) <= not(layer1_outputs(6586));
    layer2_outputs(7337) <= not(layer1_outputs(5228)) or (layer1_outputs(3899));
    layer2_outputs(7338) <= not((layer1_outputs(5852)) xor (layer1_outputs(6371)));
    layer2_outputs(7339) <= '0';
    layer2_outputs(7340) <= not(layer1_outputs(5603)) or (layer1_outputs(9913));
    layer2_outputs(7341) <= not((layer1_outputs(6668)) or (layer1_outputs(7002)));
    layer2_outputs(7342) <= (layer1_outputs(2195)) and (layer1_outputs(1459));
    layer2_outputs(7343) <= not((layer1_outputs(5361)) or (layer1_outputs(2197)));
    layer2_outputs(7344) <= layer1_outputs(692);
    layer2_outputs(7345) <= (layer1_outputs(9484)) or (layer1_outputs(7100));
    layer2_outputs(7346) <= (layer1_outputs(5962)) and not (layer1_outputs(5398));
    layer2_outputs(7347) <= not(layer1_outputs(7202)) or (layer1_outputs(144));
    layer2_outputs(7348) <= (layer1_outputs(1348)) or (layer1_outputs(9172));
    layer2_outputs(7349) <= not(layer1_outputs(680));
    layer2_outputs(7350) <= (layer1_outputs(5762)) and not (layer1_outputs(487));
    layer2_outputs(7351) <= not(layer1_outputs(2761));
    layer2_outputs(7352) <= (layer1_outputs(2406)) and not (layer1_outputs(7135));
    layer2_outputs(7353) <= not(layer1_outputs(5874));
    layer2_outputs(7354) <= layer1_outputs(3836);
    layer2_outputs(7355) <= layer1_outputs(2453);
    layer2_outputs(7356) <= not((layer1_outputs(4512)) xor (layer1_outputs(1426)));
    layer2_outputs(7357) <= (layer1_outputs(2808)) and not (layer1_outputs(7223));
    layer2_outputs(7358) <= not(layer1_outputs(9236));
    layer2_outputs(7359) <= not((layer1_outputs(5919)) or (layer1_outputs(2640)));
    layer2_outputs(7360) <= not(layer1_outputs(9422)) or (layer1_outputs(3308));
    layer2_outputs(7361) <= not(layer1_outputs(3768)) or (layer1_outputs(3333));
    layer2_outputs(7362) <= not(layer1_outputs(6331));
    layer2_outputs(7363) <= not(layer1_outputs(9370));
    layer2_outputs(7364) <= not(layer1_outputs(2244)) or (layer1_outputs(5123));
    layer2_outputs(7365) <= (layer1_outputs(137)) and not (layer1_outputs(6959));
    layer2_outputs(7366) <= layer1_outputs(2134);
    layer2_outputs(7367) <= layer1_outputs(3956);
    layer2_outputs(7368) <= not((layer1_outputs(3055)) xor (layer1_outputs(9960)));
    layer2_outputs(7369) <= layer1_outputs(4102);
    layer2_outputs(7370) <= not((layer1_outputs(2915)) or (layer1_outputs(7221)));
    layer2_outputs(7371) <= (layer1_outputs(6493)) and (layer1_outputs(4289));
    layer2_outputs(7372) <= layer1_outputs(2822);
    layer2_outputs(7373) <= layer1_outputs(4397);
    layer2_outputs(7374) <= (layer1_outputs(2576)) and not (layer1_outputs(1803));
    layer2_outputs(7375) <= not(layer1_outputs(2954));
    layer2_outputs(7376) <= not(layer1_outputs(9945));
    layer2_outputs(7377) <= layer1_outputs(2095);
    layer2_outputs(7378) <= not(layer1_outputs(392));
    layer2_outputs(7379) <= not((layer1_outputs(3511)) or (layer1_outputs(8185)));
    layer2_outputs(7380) <= not(layer1_outputs(3009));
    layer2_outputs(7381) <= (layer1_outputs(4420)) or (layer1_outputs(9588));
    layer2_outputs(7382) <= layer1_outputs(9600);
    layer2_outputs(7383) <= not(layer1_outputs(7000));
    layer2_outputs(7384) <= (layer1_outputs(4248)) and not (layer1_outputs(6082));
    layer2_outputs(7385) <= layer1_outputs(2933);
    layer2_outputs(7386) <= layer1_outputs(4029);
    layer2_outputs(7387) <= layer1_outputs(5161);
    layer2_outputs(7388) <= not(layer1_outputs(6603));
    layer2_outputs(7389) <= not(layer1_outputs(1164));
    layer2_outputs(7390) <= (layer1_outputs(3974)) and (layer1_outputs(5958));
    layer2_outputs(7391) <= not(layer1_outputs(8826)) or (layer1_outputs(9109));
    layer2_outputs(7392) <= not(layer1_outputs(1795));
    layer2_outputs(7393) <= not(layer1_outputs(1153)) or (layer1_outputs(4362));
    layer2_outputs(7394) <= not(layer1_outputs(1625)) or (layer1_outputs(4525));
    layer2_outputs(7395) <= layer1_outputs(2295);
    layer2_outputs(7396) <= layer1_outputs(6262);
    layer2_outputs(7397) <= layer1_outputs(6716);
    layer2_outputs(7398) <= not((layer1_outputs(9173)) and (layer1_outputs(4004)));
    layer2_outputs(7399) <= (layer1_outputs(416)) or (layer1_outputs(10155));
    layer2_outputs(7400) <= (layer1_outputs(4878)) or (layer1_outputs(8119));
    layer2_outputs(7401) <= (layer1_outputs(127)) and not (layer1_outputs(7024));
    layer2_outputs(7402) <= not(layer1_outputs(7004)) or (layer1_outputs(3297));
    layer2_outputs(7403) <= not(layer1_outputs(3933)) or (layer1_outputs(9255));
    layer2_outputs(7404) <= layer1_outputs(427);
    layer2_outputs(7405) <= layer1_outputs(5849);
    layer2_outputs(7406) <= not(layer1_outputs(4616));
    layer2_outputs(7407) <= not(layer1_outputs(6784));
    layer2_outputs(7408) <= (layer1_outputs(7486)) or (layer1_outputs(494));
    layer2_outputs(7409) <= layer1_outputs(7085);
    layer2_outputs(7410) <= not(layer1_outputs(4557));
    layer2_outputs(7411) <= not(layer1_outputs(6661));
    layer2_outputs(7412) <= not(layer1_outputs(5892));
    layer2_outputs(7413) <= layer1_outputs(5528);
    layer2_outputs(7414) <= not(layer1_outputs(2592));
    layer2_outputs(7415) <= (layer1_outputs(1669)) and not (layer1_outputs(5415));
    layer2_outputs(7416) <= not(layer1_outputs(8811));
    layer2_outputs(7417) <= not(layer1_outputs(7823));
    layer2_outputs(7418) <= not((layer1_outputs(10087)) or (layer1_outputs(8012)));
    layer2_outputs(7419) <= not(layer1_outputs(9976));
    layer2_outputs(7420) <= layer1_outputs(4326);
    layer2_outputs(7421) <= layer1_outputs(9713);
    layer2_outputs(7422) <= layer1_outputs(8702);
    layer2_outputs(7423) <= not((layer1_outputs(1564)) and (layer1_outputs(3525)));
    layer2_outputs(7424) <= not(layer1_outputs(3354));
    layer2_outputs(7425) <= not((layer1_outputs(6492)) xor (layer1_outputs(5221)));
    layer2_outputs(7426) <= not(layer1_outputs(2140)) or (layer1_outputs(6690));
    layer2_outputs(7427) <= not(layer1_outputs(7761));
    layer2_outputs(7428) <= (layer1_outputs(7069)) or (layer1_outputs(5325));
    layer2_outputs(7429) <= not(layer1_outputs(10091));
    layer2_outputs(7430) <= (layer1_outputs(8192)) and not (layer1_outputs(530));
    layer2_outputs(7431) <= (layer1_outputs(3477)) and not (layer1_outputs(7504));
    layer2_outputs(7432) <= layer1_outputs(2317);
    layer2_outputs(7433) <= not(layer1_outputs(7891));
    layer2_outputs(7434) <= (layer1_outputs(5369)) and not (layer1_outputs(7166));
    layer2_outputs(7435) <= layer1_outputs(5040);
    layer2_outputs(7436) <= (layer1_outputs(1473)) and (layer1_outputs(5473));
    layer2_outputs(7437) <= not((layer1_outputs(1408)) xor (layer1_outputs(6373)));
    layer2_outputs(7438) <= not(layer1_outputs(6190)) or (layer1_outputs(9664));
    layer2_outputs(7439) <= not(layer1_outputs(4250));
    layer2_outputs(7440) <= (layer1_outputs(9951)) or (layer1_outputs(1875));
    layer2_outputs(7441) <= layer1_outputs(8991);
    layer2_outputs(7442) <= layer1_outputs(3531);
    layer2_outputs(7443) <= (layer1_outputs(5116)) or (layer1_outputs(4292));
    layer2_outputs(7444) <= (layer1_outputs(2770)) and (layer1_outputs(7551));
    layer2_outputs(7445) <= not(layer1_outputs(9910));
    layer2_outputs(7446) <= '0';
    layer2_outputs(7447) <= (layer1_outputs(9613)) and (layer1_outputs(1780));
    layer2_outputs(7448) <= (layer1_outputs(2670)) or (layer1_outputs(7754));
    layer2_outputs(7449) <= layer1_outputs(2810);
    layer2_outputs(7450) <= (layer1_outputs(650)) or (layer1_outputs(3988));
    layer2_outputs(7451) <= not(layer1_outputs(5806)) or (layer1_outputs(1410));
    layer2_outputs(7452) <= not(layer1_outputs(5576));
    layer2_outputs(7453) <= not(layer1_outputs(2681));
    layer2_outputs(7454) <= (layer1_outputs(6843)) xor (layer1_outputs(4098));
    layer2_outputs(7455) <= layer1_outputs(9916);
    layer2_outputs(7456) <= layer1_outputs(2608);
    layer2_outputs(7457) <= (layer1_outputs(7703)) xor (layer1_outputs(3709));
    layer2_outputs(7458) <= not(layer1_outputs(222));
    layer2_outputs(7459) <= not(layer1_outputs(1892));
    layer2_outputs(7460) <= layer1_outputs(1404);
    layer2_outputs(7461) <= '0';
    layer2_outputs(7462) <= (layer1_outputs(1014)) and not (layer1_outputs(1117));
    layer2_outputs(7463) <= layer1_outputs(3157);
    layer2_outputs(7464) <= layer1_outputs(319);
    layer2_outputs(7465) <= not((layer1_outputs(3280)) xor (layer1_outputs(272)));
    layer2_outputs(7466) <= (layer1_outputs(8043)) and not (layer1_outputs(163));
    layer2_outputs(7467) <= not(layer1_outputs(3233));
    layer2_outputs(7468) <= not(layer1_outputs(8338)) or (layer1_outputs(5414));
    layer2_outputs(7469) <= not(layer1_outputs(6128)) or (layer1_outputs(8317));
    layer2_outputs(7470) <= not(layer1_outputs(726)) or (layer1_outputs(2234));
    layer2_outputs(7471) <= layer1_outputs(1482);
    layer2_outputs(7472) <= not(layer1_outputs(4456)) or (layer1_outputs(3375));
    layer2_outputs(7473) <= not(layer1_outputs(8425));
    layer2_outputs(7474) <= (layer1_outputs(247)) or (layer1_outputs(423));
    layer2_outputs(7475) <= not(layer1_outputs(3371));
    layer2_outputs(7476) <= not(layer1_outputs(1434));
    layer2_outputs(7477) <= not(layer1_outputs(4030));
    layer2_outputs(7478) <= not(layer1_outputs(4068)) or (layer1_outputs(1651));
    layer2_outputs(7479) <= not(layer1_outputs(8362));
    layer2_outputs(7480) <= not(layer1_outputs(5914));
    layer2_outputs(7481) <= (layer1_outputs(97)) and not (layer1_outputs(7123));
    layer2_outputs(7482) <= not(layer1_outputs(696));
    layer2_outputs(7483) <= not(layer1_outputs(2982));
    layer2_outputs(7484) <= (layer1_outputs(9856)) xor (layer1_outputs(9167));
    layer2_outputs(7485) <= not((layer1_outputs(7677)) or (layer1_outputs(5108)));
    layer2_outputs(7486) <= not(layer1_outputs(5677));
    layer2_outputs(7487) <= (layer1_outputs(6672)) and not (layer1_outputs(1274));
    layer2_outputs(7488) <= (layer1_outputs(2791)) and (layer1_outputs(8597));
    layer2_outputs(7489) <= not(layer1_outputs(8200)) or (layer1_outputs(9472));
    layer2_outputs(7490) <= not((layer1_outputs(2625)) xor (layer1_outputs(939)));
    layer2_outputs(7491) <= layer1_outputs(6357);
    layer2_outputs(7492) <= not(layer1_outputs(6563));
    layer2_outputs(7493) <= not((layer1_outputs(1355)) xor (layer1_outputs(214)));
    layer2_outputs(7494) <= '1';
    layer2_outputs(7495) <= not(layer1_outputs(9968));
    layer2_outputs(7496) <= (layer1_outputs(7738)) or (layer1_outputs(5935));
    layer2_outputs(7497) <= layer1_outputs(8412);
    layer2_outputs(7498) <= layer1_outputs(9076);
    layer2_outputs(7499) <= layer1_outputs(248);
    layer2_outputs(7500) <= not(layer1_outputs(3085)) or (layer1_outputs(71));
    layer2_outputs(7501) <= layer1_outputs(6326);
    layer2_outputs(7502) <= not(layer1_outputs(6946));
    layer2_outputs(7503) <= not(layer1_outputs(2755));
    layer2_outputs(7504) <= (layer1_outputs(6483)) and (layer1_outputs(6279));
    layer2_outputs(7505) <= layer1_outputs(6947);
    layer2_outputs(7506) <= not(layer1_outputs(10199));
    layer2_outputs(7507) <= not(layer1_outputs(2778));
    layer2_outputs(7508) <= not((layer1_outputs(3603)) or (layer1_outputs(5077)));
    layer2_outputs(7509) <= layer1_outputs(4852);
    layer2_outputs(7510) <= layer1_outputs(6289);
    layer2_outputs(7511) <= layer1_outputs(3202);
    layer2_outputs(7512) <= not((layer1_outputs(4306)) xor (layer1_outputs(7588)));
    layer2_outputs(7513) <= (layer1_outputs(6440)) and not (layer1_outputs(2414));
    layer2_outputs(7514) <= (layer1_outputs(475)) and not (layer1_outputs(9994));
    layer2_outputs(7515) <= (layer1_outputs(2368)) and not (layer1_outputs(7606));
    layer2_outputs(7516) <= not(layer1_outputs(3365));
    layer2_outputs(7517) <= not((layer1_outputs(4170)) xor (layer1_outputs(9784)));
    layer2_outputs(7518) <= not((layer1_outputs(3815)) xor (layer1_outputs(1597)));
    layer2_outputs(7519) <= (layer1_outputs(9220)) and not (layer1_outputs(6791));
    layer2_outputs(7520) <= not(layer1_outputs(7061));
    layer2_outputs(7521) <= not((layer1_outputs(3977)) or (layer1_outputs(5103)));
    layer2_outputs(7522) <= not(layer1_outputs(3177));
    layer2_outputs(7523) <= not((layer1_outputs(6772)) xor (layer1_outputs(3734)));
    layer2_outputs(7524) <= not((layer1_outputs(4075)) and (layer1_outputs(2282)));
    layer2_outputs(7525) <= layer1_outputs(3846);
    layer2_outputs(7526) <= layer1_outputs(2750);
    layer2_outputs(7527) <= not((layer1_outputs(10228)) and (layer1_outputs(9639)));
    layer2_outputs(7528) <= layer1_outputs(10025);
    layer2_outputs(7529) <= not(layer1_outputs(8558));
    layer2_outputs(7530) <= not((layer1_outputs(75)) xor (layer1_outputs(9198)));
    layer2_outputs(7531) <= (layer1_outputs(4279)) xor (layer1_outputs(6386));
    layer2_outputs(7532) <= (layer1_outputs(1382)) xor (layer1_outputs(3388));
    layer2_outputs(7533) <= (layer1_outputs(2193)) and not (layer1_outputs(1652));
    layer2_outputs(7534) <= layer1_outputs(6161);
    layer2_outputs(7535) <= (layer1_outputs(1267)) and not (layer1_outputs(6827));
    layer2_outputs(7536) <= not(layer1_outputs(4352));
    layer2_outputs(7537) <= '0';
    layer2_outputs(7538) <= not((layer1_outputs(8577)) or (layer1_outputs(1061)));
    layer2_outputs(7539) <= (layer1_outputs(4226)) or (layer1_outputs(3567));
    layer2_outputs(7540) <= not(layer1_outputs(7679));
    layer2_outputs(7541) <= (layer1_outputs(3623)) and (layer1_outputs(7375));
    layer2_outputs(7542) <= layer1_outputs(5559);
    layer2_outputs(7543) <= not(layer1_outputs(5891));
    layer2_outputs(7544) <= not(layer1_outputs(2122));
    layer2_outputs(7545) <= layer1_outputs(7249);
    layer2_outputs(7546) <= not(layer1_outputs(955));
    layer2_outputs(7547) <= (layer1_outputs(6698)) and not (layer1_outputs(3322));
    layer2_outputs(7548) <= layer1_outputs(2094);
    layer2_outputs(7549) <= not((layer1_outputs(7586)) or (layer1_outputs(7987)));
    layer2_outputs(7550) <= not((layer1_outputs(9839)) xor (layer1_outputs(9413)));
    layer2_outputs(7551) <= not((layer1_outputs(6927)) xor (layer1_outputs(7889)));
    layer2_outputs(7552) <= not(layer1_outputs(9891));
    layer2_outputs(7553) <= not(layer1_outputs(5640)) or (layer1_outputs(9022));
    layer2_outputs(7554) <= not(layer1_outputs(6378));
    layer2_outputs(7555) <= (layer1_outputs(1847)) and not (layer1_outputs(6797));
    layer2_outputs(7556) <= (layer1_outputs(2207)) and not (layer1_outputs(3319));
    layer2_outputs(7557) <= not((layer1_outputs(3009)) xor (layer1_outputs(39)));
    layer2_outputs(7558) <= (layer1_outputs(5514)) xor (layer1_outputs(2538));
    layer2_outputs(7559) <= not(layer1_outputs(2)) or (layer1_outputs(2604));
    layer2_outputs(7560) <= layer1_outputs(1502);
    layer2_outputs(7561) <= layer1_outputs(9930);
    layer2_outputs(7562) <= not(layer1_outputs(9961));
    layer2_outputs(7563) <= not((layer1_outputs(7956)) xor (layer1_outputs(4161)));
    layer2_outputs(7564) <= layer1_outputs(2533);
    layer2_outputs(7565) <= (layer1_outputs(10163)) or (layer1_outputs(6844));
    layer2_outputs(7566) <= not((layer1_outputs(10138)) or (layer1_outputs(8160)));
    layer2_outputs(7567) <= layer1_outputs(3455);
    layer2_outputs(7568) <= not(layer1_outputs(1982));
    layer2_outputs(7569) <= not((layer1_outputs(7807)) and (layer1_outputs(4910)));
    layer2_outputs(7570) <= layer1_outputs(5049);
    layer2_outputs(7571) <= (layer1_outputs(122)) and (layer1_outputs(4798));
    layer2_outputs(7572) <= not(layer1_outputs(9988));
    layer2_outputs(7573) <= not((layer1_outputs(1822)) xor (layer1_outputs(7125)));
    layer2_outputs(7574) <= not(layer1_outputs(3967)) or (layer1_outputs(591));
    layer2_outputs(7575) <= '1';
    layer2_outputs(7576) <= layer1_outputs(5421);
    layer2_outputs(7577) <= (layer1_outputs(5241)) and not (layer1_outputs(7844));
    layer2_outputs(7578) <= not((layer1_outputs(4844)) xor (layer1_outputs(9335)));
    layer2_outputs(7579) <= not(layer1_outputs(6276));
    layer2_outputs(7580) <= not(layer1_outputs(9563));
    layer2_outputs(7581) <= not(layer1_outputs(5005)) or (layer1_outputs(8356));
    layer2_outputs(7582) <= (layer1_outputs(7839)) and not (layer1_outputs(4846));
    layer2_outputs(7583) <= not(layer1_outputs(5574)) or (layer1_outputs(752));
    layer2_outputs(7584) <= not((layer1_outputs(1762)) and (layer1_outputs(7222)));
    layer2_outputs(7585) <= (layer1_outputs(9898)) xor (layer1_outputs(4972));
    layer2_outputs(7586) <= '0';
    layer2_outputs(7587) <= not(layer1_outputs(6677));
    layer2_outputs(7588) <= not((layer1_outputs(3569)) xor (layer1_outputs(9744)));
    layer2_outputs(7589) <= not((layer1_outputs(5994)) or (layer1_outputs(6824)));
    layer2_outputs(7590) <= layer1_outputs(6265);
    layer2_outputs(7591) <= not((layer1_outputs(8445)) xor (layer1_outputs(4806)));
    layer2_outputs(7592) <= not(layer1_outputs(393)) or (layer1_outputs(9345));
    layer2_outputs(7593) <= layer1_outputs(549);
    layer2_outputs(7594) <= not(layer1_outputs(243));
    layer2_outputs(7595) <= (layer1_outputs(2267)) and not (layer1_outputs(4824));
    layer2_outputs(7596) <= not(layer1_outputs(6547));
    layer2_outputs(7597) <= (layer1_outputs(7686)) xor (layer1_outputs(1820));
    layer2_outputs(7598) <= not(layer1_outputs(957)) or (layer1_outputs(3652));
    layer2_outputs(7599) <= not(layer1_outputs(8687));
    layer2_outputs(7600) <= not((layer1_outputs(3083)) xor (layer1_outputs(9808)));
    layer2_outputs(7601) <= not(layer1_outputs(887));
    layer2_outputs(7602) <= not(layer1_outputs(3078));
    layer2_outputs(7603) <= not((layer1_outputs(2664)) xor (layer1_outputs(6249)));
    layer2_outputs(7604) <= layer1_outputs(5391);
    layer2_outputs(7605) <= not(layer1_outputs(3523)) or (layer1_outputs(1118));
    layer2_outputs(7606) <= not(layer1_outputs(438));
    layer2_outputs(7607) <= (layer1_outputs(399)) or (layer1_outputs(5437));
    layer2_outputs(7608) <= (layer1_outputs(3267)) and not (layer1_outputs(8958));
    layer2_outputs(7609) <= layer1_outputs(5828);
    layer2_outputs(7610) <= not((layer1_outputs(5443)) and (layer1_outputs(1391)));
    layer2_outputs(7611) <= not(layer1_outputs(9596));
    layer2_outputs(7612) <= not(layer1_outputs(2788));
    layer2_outputs(7613) <= not(layer1_outputs(2996)) or (layer1_outputs(1920));
    layer2_outputs(7614) <= not((layer1_outputs(3185)) or (layer1_outputs(9838)));
    layer2_outputs(7615) <= layer1_outputs(4340);
    layer2_outputs(7616) <= layer1_outputs(7049);
    layer2_outputs(7617) <= layer1_outputs(7686);
    layer2_outputs(7618) <= (layer1_outputs(8752)) xor (layer1_outputs(8917));
    layer2_outputs(7619) <= (layer1_outputs(4262)) xor (layer1_outputs(4853));
    layer2_outputs(7620) <= not((layer1_outputs(9132)) and (layer1_outputs(8281)));
    layer2_outputs(7621) <= not(layer1_outputs(9511));
    layer2_outputs(7622) <= not(layer1_outputs(7239));
    layer2_outputs(7623) <= (layer1_outputs(6342)) xor (layer1_outputs(3670));
    layer2_outputs(7624) <= layer1_outputs(8901);
    layer2_outputs(7625) <= (layer1_outputs(9924)) xor (layer1_outputs(8107));
    layer2_outputs(7626) <= not(layer1_outputs(9678));
    layer2_outputs(7627) <= not(layer1_outputs(9244)) or (layer1_outputs(3200));
    layer2_outputs(7628) <= layer1_outputs(2787);
    layer2_outputs(7629) <= not(layer1_outputs(4950));
    layer2_outputs(7630) <= not((layer1_outputs(9521)) and (layer1_outputs(3350)));
    layer2_outputs(7631) <= (layer1_outputs(10189)) and (layer1_outputs(1267));
    layer2_outputs(7632) <= layer1_outputs(7165);
    layer2_outputs(7633) <= not(layer1_outputs(5881));
    layer2_outputs(7634) <= layer1_outputs(643);
    layer2_outputs(7635) <= not(layer1_outputs(2297)) or (layer1_outputs(8841));
    layer2_outputs(7636) <= not(layer1_outputs(4095));
    layer2_outputs(7637) <= not(layer1_outputs(4591)) or (layer1_outputs(5650));
    layer2_outputs(7638) <= (layer1_outputs(9243)) and not (layer1_outputs(2886));
    layer2_outputs(7639) <= (layer1_outputs(5820)) and not (layer1_outputs(4879));
    layer2_outputs(7640) <= layer1_outputs(5149);
    layer2_outputs(7641) <= layer1_outputs(4788);
    layer2_outputs(7642) <= layer1_outputs(2485);
    layer2_outputs(7643) <= not(layer1_outputs(7184)) or (layer1_outputs(9328));
    layer2_outputs(7644) <= not(layer1_outputs(3915));
    layer2_outputs(7645) <= layer1_outputs(6935);
    layer2_outputs(7646) <= layer1_outputs(6863);
    layer2_outputs(7647) <= (layer1_outputs(10004)) and not (layer1_outputs(524));
    layer2_outputs(7648) <= not((layer1_outputs(5332)) and (layer1_outputs(6287)));
    layer2_outputs(7649) <= (layer1_outputs(9895)) and not (layer1_outputs(1503));
    layer2_outputs(7650) <= layer1_outputs(4846);
    layer2_outputs(7651) <= not((layer1_outputs(1520)) or (layer1_outputs(1815)));
    layer2_outputs(7652) <= not(layer1_outputs(5955));
    layer2_outputs(7653) <= layer1_outputs(5179);
    layer2_outputs(7654) <= (layer1_outputs(413)) or (layer1_outputs(2730));
    layer2_outputs(7655) <= (layer1_outputs(3421)) xor (layer1_outputs(4698));
    layer2_outputs(7656) <= not((layer1_outputs(5355)) or (layer1_outputs(3369)));
    layer2_outputs(7657) <= (layer1_outputs(6269)) or (layer1_outputs(2790));
    layer2_outputs(7658) <= not(layer1_outputs(1232));
    layer2_outputs(7659) <= layer1_outputs(9404);
    layer2_outputs(7660) <= not((layer1_outputs(5817)) and (layer1_outputs(1133)));
    layer2_outputs(7661) <= layer1_outputs(1847);
    layer2_outputs(7662) <= (layer1_outputs(1251)) or (layer1_outputs(5890));
    layer2_outputs(7663) <= not((layer1_outputs(8343)) or (layer1_outputs(349)));
    layer2_outputs(7664) <= not(layer1_outputs(4050));
    layer2_outputs(7665) <= (layer1_outputs(3775)) and not (layer1_outputs(6850));
    layer2_outputs(7666) <= (layer1_outputs(5023)) and not (layer1_outputs(10046));
    layer2_outputs(7667) <= (layer1_outputs(5196)) and not (layer1_outputs(1901));
    layer2_outputs(7668) <= not(layer1_outputs(9626));
    layer2_outputs(7669) <= layer1_outputs(1071);
    layer2_outputs(7670) <= (layer1_outputs(2902)) xor (layer1_outputs(3881));
    layer2_outputs(7671) <= (layer1_outputs(7861)) or (layer1_outputs(10063));
    layer2_outputs(7672) <= (layer1_outputs(7400)) and not (layer1_outputs(1405));
    layer2_outputs(7673) <= layer1_outputs(8960);
    layer2_outputs(7674) <= not((layer1_outputs(3883)) and (layer1_outputs(1545)));
    layer2_outputs(7675) <= layer1_outputs(8886);
    layer2_outputs(7676) <= layer1_outputs(2615);
    layer2_outputs(7677) <= not((layer1_outputs(7639)) or (layer1_outputs(5228)));
    layer2_outputs(7678) <= not(layer1_outputs(1326)) or (layer1_outputs(7359));
    layer2_outputs(7679) <= not(layer1_outputs(4163));
    layer2_outputs(7680) <= layer1_outputs(9681);
    layer2_outputs(7681) <= not(layer1_outputs(2482)) or (layer1_outputs(9382));
    layer2_outputs(7682) <= not(layer1_outputs(688)) or (layer1_outputs(5540));
    layer2_outputs(7683) <= layer1_outputs(8551);
    layer2_outputs(7684) <= layer1_outputs(6496);
    layer2_outputs(7685) <= layer1_outputs(7972);
    layer2_outputs(7686) <= not(layer1_outputs(6554));
    layer2_outputs(7687) <= (layer1_outputs(4778)) and not (layer1_outputs(1026));
    layer2_outputs(7688) <= layer1_outputs(7813);
    layer2_outputs(7689) <= layer1_outputs(1062);
    layer2_outputs(7690) <= (layer1_outputs(956)) xor (layer1_outputs(9671));
    layer2_outputs(7691) <= not((layer1_outputs(2023)) xor (layer1_outputs(4119)));
    layer2_outputs(7692) <= (layer1_outputs(866)) xor (layer1_outputs(5232));
    layer2_outputs(7693) <= not((layer1_outputs(5950)) xor (layer1_outputs(104)));
    layer2_outputs(7694) <= not((layer1_outputs(103)) or (layer1_outputs(9066)));
    layer2_outputs(7695) <= (layer1_outputs(102)) and (layer1_outputs(6445));
    layer2_outputs(7696) <= (layer1_outputs(1295)) xor (layer1_outputs(2931));
    layer2_outputs(7697) <= not(layer1_outputs(3933)) or (layer1_outputs(6105));
    layer2_outputs(7698) <= (layer1_outputs(2932)) xor (layer1_outputs(9368));
    layer2_outputs(7699) <= not((layer1_outputs(7798)) and (layer1_outputs(7447)));
    layer2_outputs(7700) <= not((layer1_outputs(1784)) and (layer1_outputs(9819)));
    layer2_outputs(7701) <= not(layer1_outputs(8190));
    layer2_outputs(7702) <= (layer1_outputs(3931)) and not (layer1_outputs(6498));
    layer2_outputs(7703) <= layer1_outputs(9350);
    layer2_outputs(7704) <= (layer1_outputs(5006)) and not (layer1_outputs(8859));
    layer2_outputs(7705) <= (layer1_outputs(9841)) and (layer1_outputs(6344));
    layer2_outputs(7706) <= not(layer1_outputs(6951));
    layer2_outputs(7707) <= (layer1_outputs(3014)) or (layer1_outputs(3860));
    layer2_outputs(7708) <= layer1_outputs(115);
    layer2_outputs(7709) <= layer1_outputs(3596);
    layer2_outputs(7710) <= not(layer1_outputs(6935)) or (layer1_outputs(4499));
    layer2_outputs(7711) <= layer1_outputs(9764);
    layer2_outputs(7712) <= not(layer1_outputs(10230));
    layer2_outputs(7713) <= not((layer1_outputs(898)) and (layer1_outputs(7608)));
    layer2_outputs(7714) <= (layer1_outputs(6945)) and not (layer1_outputs(7243));
    layer2_outputs(7715) <= not(layer1_outputs(9155)) or (layer1_outputs(4505));
    layer2_outputs(7716) <= not(layer1_outputs(10210));
    layer2_outputs(7717) <= not(layer1_outputs(1393));
    layer2_outputs(7718) <= (layer1_outputs(8252)) and (layer1_outputs(2033));
    layer2_outputs(7719) <= not(layer1_outputs(949));
    layer2_outputs(7720) <= (layer1_outputs(2722)) xor (layer1_outputs(9620));
    layer2_outputs(7721) <= not(layer1_outputs(5566)) or (layer1_outputs(1077));
    layer2_outputs(7722) <= not(layer1_outputs(1808));
    layer2_outputs(7723) <= (layer1_outputs(6324)) and (layer1_outputs(5469));
    layer2_outputs(7724) <= not(layer1_outputs(6507));
    layer2_outputs(7725) <= (layer1_outputs(5444)) and not (layer1_outputs(1032));
    layer2_outputs(7726) <= not(layer1_outputs(8313));
    layer2_outputs(7727) <= layer1_outputs(6141);
    layer2_outputs(7728) <= not(layer1_outputs(4546));
    layer2_outputs(7729) <= (layer1_outputs(534)) and not (layer1_outputs(1553));
    layer2_outputs(7730) <= (layer1_outputs(376)) and not (layer1_outputs(4734));
    layer2_outputs(7731) <= not((layer1_outputs(8278)) or (layer1_outputs(979)));
    layer2_outputs(7732) <= (layer1_outputs(155)) and not (layer1_outputs(4458));
    layer2_outputs(7733) <= (layer1_outputs(2738)) or (layer1_outputs(8954));
    layer2_outputs(7734) <= not(layer1_outputs(677));
    layer2_outputs(7735) <= not(layer1_outputs(5860)) or (layer1_outputs(8387));
    layer2_outputs(7736) <= not(layer1_outputs(8066)) or (layer1_outputs(70));
    layer2_outputs(7737) <= not(layer1_outputs(1097));
    layer2_outputs(7738) <= not((layer1_outputs(3875)) or (layer1_outputs(4343)));
    layer2_outputs(7739) <= not((layer1_outputs(4294)) and (layer1_outputs(5773)));
    layer2_outputs(7740) <= not(layer1_outputs(5408));
    layer2_outputs(7741) <= not(layer1_outputs(5792));
    layer2_outputs(7742) <= layer1_outputs(2002);
    layer2_outputs(7743) <= not((layer1_outputs(22)) and (layer1_outputs(8228)));
    layer2_outputs(7744) <= not(layer1_outputs(8165)) or (layer1_outputs(6372));
    layer2_outputs(7745) <= layer1_outputs(8110);
    layer2_outputs(7746) <= not(layer1_outputs(5165));
    layer2_outputs(7747) <= layer1_outputs(9182);
    layer2_outputs(7748) <= not(layer1_outputs(7952)) or (layer1_outputs(7124));
    layer2_outputs(7749) <= not(layer1_outputs(6113)) or (layer1_outputs(4370));
    layer2_outputs(7750) <= not(layer1_outputs(5572));
    layer2_outputs(7751) <= not((layer1_outputs(6202)) xor (layer1_outputs(3935)));
    layer2_outputs(7752) <= (layer1_outputs(9912)) xor (layer1_outputs(3785));
    layer2_outputs(7753) <= layer1_outputs(7675);
    layer2_outputs(7754) <= '0';
    layer2_outputs(7755) <= not(layer1_outputs(8988));
    layer2_outputs(7756) <= (layer1_outputs(6584)) or (layer1_outputs(250));
    layer2_outputs(7757) <= layer1_outputs(8529);
    layer2_outputs(7758) <= layer1_outputs(7875);
    layer2_outputs(7759) <= (layer1_outputs(9975)) and (layer1_outputs(8819));
    layer2_outputs(7760) <= not(layer1_outputs(4651));
    layer2_outputs(7761) <= not((layer1_outputs(871)) or (layer1_outputs(1462)));
    layer2_outputs(7762) <= not(layer1_outputs(8657));
    layer2_outputs(7763) <= layer1_outputs(7656);
    layer2_outputs(7764) <= layer1_outputs(6181);
    layer2_outputs(7765) <= layer1_outputs(5124);
    layer2_outputs(7766) <= layer1_outputs(9937);
    layer2_outputs(7767) <= not((layer1_outputs(1553)) and (layer1_outputs(4015)));
    layer2_outputs(7768) <= not(layer1_outputs(8505));
    layer2_outputs(7769) <= layer1_outputs(3909);
    layer2_outputs(7770) <= (layer1_outputs(4349)) and not (layer1_outputs(576));
    layer2_outputs(7771) <= layer1_outputs(5109);
    layer2_outputs(7772) <= (layer1_outputs(1656)) xor (layer1_outputs(4750));
    layer2_outputs(7773) <= not(layer1_outputs(4713));
    layer2_outputs(7774) <= (layer1_outputs(6549)) and not (layer1_outputs(4550));
    layer2_outputs(7775) <= layer1_outputs(3759);
    layer2_outputs(7776) <= not((layer1_outputs(6185)) or (layer1_outputs(5707)));
    layer2_outputs(7777) <= (layer1_outputs(3884)) and (layer1_outputs(4243));
    layer2_outputs(7778) <= (layer1_outputs(9559)) or (layer1_outputs(4199));
    layer2_outputs(7779) <= (layer1_outputs(8301)) xor (layer1_outputs(2562));
    layer2_outputs(7780) <= layer1_outputs(2233);
    layer2_outputs(7781) <= '0';
    layer2_outputs(7782) <= layer1_outputs(8711);
    layer2_outputs(7783) <= not((layer1_outputs(7759)) or (layer1_outputs(3431)));
    layer2_outputs(7784) <= (layer1_outputs(5386)) xor (layer1_outputs(1194));
    layer2_outputs(7785) <= not((layer1_outputs(7080)) xor (layer1_outputs(7249)));
    layer2_outputs(7786) <= not((layer1_outputs(3328)) and (layer1_outputs(2285)));
    layer2_outputs(7787) <= layer1_outputs(6083);
    layer2_outputs(7788) <= not(layer1_outputs(5028));
    layer2_outputs(7789) <= layer1_outputs(6864);
    layer2_outputs(7790) <= not((layer1_outputs(2649)) xor (layer1_outputs(1192)));
    layer2_outputs(7791) <= not((layer1_outputs(7138)) and (layer1_outputs(6189)));
    layer2_outputs(7792) <= not((layer1_outputs(5363)) xor (layer1_outputs(9241)));
    layer2_outputs(7793) <= layer1_outputs(3224);
    layer2_outputs(7794) <= not(layer1_outputs(3508));
    layer2_outputs(7795) <= not(layer1_outputs(8130)) or (layer1_outputs(3566));
    layer2_outputs(7796) <= (layer1_outputs(2701)) and not (layer1_outputs(3400));
    layer2_outputs(7797) <= layer1_outputs(5059);
    layer2_outputs(7798) <= not((layer1_outputs(3058)) or (layer1_outputs(7143)));
    layer2_outputs(7799) <= '0';
    layer2_outputs(7800) <= layer1_outputs(4954);
    layer2_outputs(7801) <= not(layer1_outputs(7523)) or (layer1_outputs(7544));
    layer2_outputs(7802) <= (layer1_outputs(8986)) and (layer1_outputs(6829));
    layer2_outputs(7803) <= not(layer1_outputs(8512)) or (layer1_outputs(5427));
    layer2_outputs(7804) <= not(layer1_outputs(2531));
    layer2_outputs(7805) <= not(layer1_outputs(5404));
    layer2_outputs(7806) <= (layer1_outputs(8167)) xor (layer1_outputs(1309));
    layer2_outputs(7807) <= (layer1_outputs(802)) or (layer1_outputs(4159));
    layer2_outputs(7808) <= layer1_outputs(2801);
    layer2_outputs(7809) <= not((layer1_outputs(1115)) and (layer1_outputs(6803)));
    layer2_outputs(7810) <= layer1_outputs(3034);
    layer2_outputs(7811) <= layer1_outputs(7500);
    layer2_outputs(7812) <= not(layer1_outputs(8976)) or (layer1_outputs(2631));
    layer2_outputs(7813) <= not(layer1_outputs(2220)) or (layer1_outputs(7966));
    layer2_outputs(7814) <= not((layer1_outputs(4076)) and (layer1_outputs(1021)));
    layer2_outputs(7815) <= (layer1_outputs(9885)) and not (layer1_outputs(4913));
    layer2_outputs(7816) <= (layer1_outputs(6686)) and (layer1_outputs(835));
    layer2_outputs(7817) <= not(layer1_outputs(324));
    layer2_outputs(7818) <= not((layer1_outputs(5901)) xor (layer1_outputs(1542)));
    layer2_outputs(7819) <= not(layer1_outputs(6024)) or (layer1_outputs(3262));
    layer2_outputs(7820) <= layer1_outputs(4357);
    layer2_outputs(7821) <= (layer1_outputs(7740)) and not (layer1_outputs(2930));
    layer2_outputs(7822) <= not(layer1_outputs(4491)) or (layer1_outputs(876));
    layer2_outputs(7823) <= layer1_outputs(3502);
    layer2_outputs(7824) <= not(layer1_outputs(5656)) or (layer1_outputs(8754));
    layer2_outputs(7825) <= (layer1_outputs(1347)) xor (layer1_outputs(9775));
    layer2_outputs(7826) <= (layer1_outputs(6849)) xor (layer1_outputs(5481));
    layer2_outputs(7827) <= layer1_outputs(333);
    layer2_outputs(7828) <= layer1_outputs(7130);
    layer2_outputs(7829) <= layer1_outputs(8391);
    layer2_outputs(7830) <= not(layer1_outputs(7437)) or (layer1_outputs(9394));
    layer2_outputs(7831) <= not((layer1_outputs(7150)) or (layer1_outputs(9477)));
    layer2_outputs(7832) <= layer1_outputs(2277);
    layer2_outputs(7833) <= (layer1_outputs(5797)) and (layer1_outputs(4818));
    layer2_outputs(7834) <= not(layer1_outputs(613)) or (layer1_outputs(583));
    layer2_outputs(7835) <= (layer1_outputs(2478)) xor (layer1_outputs(9401));
    layer2_outputs(7836) <= not(layer1_outputs(2241)) or (layer1_outputs(1360));
    layer2_outputs(7837) <= not(layer1_outputs(1677));
    layer2_outputs(7838) <= not(layer1_outputs(8475));
    layer2_outputs(7839) <= not((layer1_outputs(2997)) xor (layer1_outputs(5456)));
    layer2_outputs(7840) <= not((layer1_outputs(9233)) or (layer1_outputs(1576)));
    layer2_outputs(7841) <= layer1_outputs(7753);
    layer2_outputs(7842) <= not(layer1_outputs(9050));
    layer2_outputs(7843) <= not(layer1_outputs(3106));
    layer2_outputs(7844) <= not(layer1_outputs(6795));
    layer2_outputs(7845) <= not(layer1_outputs(9697));
    layer2_outputs(7846) <= not(layer1_outputs(7767)) or (layer1_outputs(5745));
    layer2_outputs(7847) <= layer1_outputs(862);
    layer2_outputs(7848) <= layer1_outputs(8854);
    layer2_outputs(7849) <= not(layer1_outputs(9775)) or (layer1_outputs(7005));
    layer2_outputs(7850) <= not((layer1_outputs(963)) or (layer1_outputs(2855)));
    layer2_outputs(7851) <= (layer1_outputs(1285)) or (layer1_outputs(7901));
    layer2_outputs(7852) <= layer1_outputs(7376);
    layer2_outputs(7853) <= not(layer1_outputs(4679));
    layer2_outputs(7854) <= layer1_outputs(919);
    layer2_outputs(7855) <= (layer1_outputs(5549)) and not (layer1_outputs(4285));
    layer2_outputs(7856) <= (layer1_outputs(2251)) or (layer1_outputs(6954));
    layer2_outputs(7857) <= not(layer1_outputs(4211));
    layer2_outputs(7858) <= not(layer1_outputs(2385));
    layer2_outputs(7859) <= layer1_outputs(4006);
    layer2_outputs(7860) <= not(layer1_outputs(1961));
    layer2_outputs(7861) <= not(layer1_outputs(4743));
    layer2_outputs(7862) <= not(layer1_outputs(893));
    layer2_outputs(7863) <= not((layer1_outputs(5558)) and (layer1_outputs(8319)));
    layer2_outputs(7864) <= layer1_outputs(1742);
    layer2_outputs(7865) <= not(layer1_outputs(7698));
    layer2_outputs(7866) <= not(layer1_outputs(6621));
    layer2_outputs(7867) <= not(layer1_outputs(4777)) or (layer1_outputs(4128));
    layer2_outputs(7868) <= not(layer1_outputs(827));
    layer2_outputs(7869) <= not(layer1_outputs(9470));
    layer2_outputs(7870) <= '0';
    layer2_outputs(7871) <= (layer1_outputs(9420)) and not (layer1_outputs(8839));
    layer2_outputs(7872) <= not((layer1_outputs(2988)) or (layer1_outputs(6886)));
    layer2_outputs(7873) <= not(layer1_outputs(8954)) or (layer1_outputs(6257));
    layer2_outputs(7874) <= layer1_outputs(2552);
    layer2_outputs(7875) <= not(layer1_outputs(327));
    layer2_outputs(7876) <= layer1_outputs(5199);
    layer2_outputs(7877) <= not(layer1_outputs(8696)) or (layer1_outputs(5098));
    layer2_outputs(7878) <= not((layer1_outputs(10072)) and (layer1_outputs(484)));
    layer2_outputs(7879) <= not(layer1_outputs(1074)) or (layer1_outputs(4984));
    layer2_outputs(7880) <= not(layer1_outputs(5996));
    layer2_outputs(7881) <= layer1_outputs(5734);
    layer2_outputs(7882) <= not((layer1_outputs(3051)) and (layer1_outputs(9341)));
    layer2_outputs(7883) <= not((layer1_outputs(8365)) or (layer1_outputs(7359)));
    layer2_outputs(7884) <= not(layer1_outputs(4472));
    layer2_outputs(7885) <= not(layer1_outputs(1744));
    layer2_outputs(7886) <= (layer1_outputs(6608)) or (layer1_outputs(5907));
    layer2_outputs(7887) <= layer1_outputs(4424);
    layer2_outputs(7888) <= layer1_outputs(9427);
    layer2_outputs(7889) <= layer1_outputs(6444);
    layer2_outputs(7890) <= not(layer1_outputs(83));
    layer2_outputs(7891) <= not(layer1_outputs(9861));
    layer2_outputs(7892) <= not(layer1_outputs(2780));
    layer2_outputs(7893) <= (layer1_outputs(5672)) and not (layer1_outputs(7997));
    layer2_outputs(7894) <= not(layer1_outputs(6614));
    layer2_outputs(7895) <= (layer1_outputs(2814)) and not (layer1_outputs(6936));
    layer2_outputs(7896) <= not(layer1_outputs(6695));
    layer2_outputs(7897) <= (layer1_outputs(6974)) or (layer1_outputs(9809));
    layer2_outputs(7898) <= '0';
    layer2_outputs(7899) <= not(layer1_outputs(2404));
    layer2_outputs(7900) <= (layer1_outputs(8227)) and (layer1_outputs(6979));
    layer2_outputs(7901) <= layer1_outputs(1403);
    layer2_outputs(7902) <= (layer1_outputs(6878)) and not (layer1_outputs(3145));
    layer2_outputs(7903) <= not((layer1_outputs(2263)) and (layer1_outputs(5916)));
    layer2_outputs(7904) <= not(layer1_outputs(5102));
    layer2_outputs(7905) <= not(layer1_outputs(9582)) or (layer1_outputs(1151));
    layer2_outputs(7906) <= (layer1_outputs(5833)) and not (layer1_outputs(3733));
    layer2_outputs(7907) <= not((layer1_outputs(1080)) or (layer1_outputs(1953)));
    layer2_outputs(7908) <= layer1_outputs(1255);
    layer2_outputs(7909) <= not((layer1_outputs(774)) or (layer1_outputs(1540)));
    layer2_outputs(7910) <= (layer1_outputs(9740)) and not (layer1_outputs(759));
    layer2_outputs(7911) <= layer1_outputs(2603);
    layer2_outputs(7912) <= (layer1_outputs(8409)) xor (layer1_outputs(7314));
    layer2_outputs(7913) <= not(layer1_outputs(8825));
    layer2_outputs(7914) <= not((layer1_outputs(9948)) xor (layer1_outputs(8215)));
    layer2_outputs(7915) <= not(layer1_outputs(1583));
    layer2_outputs(7916) <= not(layer1_outputs(9193)) or (layer1_outputs(665));
    layer2_outputs(7917) <= layer1_outputs(2113);
    layer2_outputs(7918) <= (layer1_outputs(3419)) and not (layer1_outputs(1567));
    layer2_outputs(7919) <= layer1_outputs(821);
    layer2_outputs(7920) <= (layer1_outputs(9425)) xor (layer1_outputs(2461));
    layer2_outputs(7921) <= not(layer1_outputs(3820));
    layer2_outputs(7922) <= not(layer1_outputs(7057)) or (layer1_outputs(150));
    layer2_outputs(7923) <= (layer1_outputs(8036)) and (layer1_outputs(1391));
    layer2_outputs(7924) <= (layer1_outputs(9363)) or (layer1_outputs(8406));
    layer2_outputs(7925) <= not(layer1_outputs(7293)) or (layer1_outputs(1285));
    layer2_outputs(7926) <= not(layer1_outputs(3604));
    layer2_outputs(7927) <= not((layer1_outputs(6088)) or (layer1_outputs(2291)));
    layer2_outputs(7928) <= (layer1_outputs(8937)) or (layer1_outputs(207));
    layer2_outputs(7929) <= (layer1_outputs(9555)) or (layer1_outputs(7848));
    layer2_outputs(7930) <= (layer1_outputs(412)) xor (layer1_outputs(7352));
    layer2_outputs(7931) <= not(layer1_outputs(2231)) or (layer1_outputs(5467));
    layer2_outputs(7932) <= not(layer1_outputs(8770));
    layer2_outputs(7933) <= layer1_outputs(7719);
    layer2_outputs(7934) <= layer1_outputs(6977);
    layer2_outputs(7935) <= not(layer1_outputs(8618)) or (layer1_outputs(3298));
    layer2_outputs(7936) <= not((layer1_outputs(6807)) and (layer1_outputs(10156)));
    layer2_outputs(7937) <= layer1_outputs(9243);
    layer2_outputs(7938) <= not(layer1_outputs(782));
    layer2_outputs(7939) <= (layer1_outputs(6879)) or (layer1_outputs(3489));
    layer2_outputs(7940) <= not(layer1_outputs(10067));
    layer2_outputs(7941) <= layer1_outputs(8936);
    layer2_outputs(7942) <= not((layer1_outputs(6974)) and (layer1_outputs(3394)));
    layer2_outputs(7943) <= not(layer1_outputs(8143));
    layer2_outputs(7944) <= layer1_outputs(404);
    layer2_outputs(7945) <= (layer1_outputs(487)) and not (layer1_outputs(184));
    layer2_outputs(7946) <= not((layer1_outputs(4418)) and (layer1_outputs(6063)));
    layer2_outputs(7947) <= not((layer1_outputs(6572)) and (layer1_outputs(7799)));
    layer2_outputs(7948) <= layer1_outputs(4593);
    layer2_outputs(7949) <= not((layer1_outputs(6305)) and (layer1_outputs(3190)));
    layer2_outputs(7950) <= not((layer1_outputs(4500)) xor (layer1_outputs(1182)));
    layer2_outputs(7951) <= (layer1_outputs(215)) and not (layer1_outputs(3512));
    layer2_outputs(7952) <= not(layer1_outputs(6940)) or (layer1_outputs(4064));
    layer2_outputs(7953) <= not(layer1_outputs(5201)) or (layer1_outputs(7550));
    layer2_outputs(7954) <= not(layer1_outputs(7061));
    layer2_outputs(7955) <= not((layer1_outputs(9703)) xor (layer1_outputs(6455)));
    layer2_outputs(7956) <= (layer1_outputs(3257)) or (layer1_outputs(9143));
    layer2_outputs(7957) <= (layer1_outputs(5310)) or (layer1_outputs(4282));
    layer2_outputs(7958) <= not(layer1_outputs(5760));
    layer2_outputs(7959) <= (layer1_outputs(5448)) or (layer1_outputs(9760));
    layer2_outputs(7960) <= not(layer1_outputs(162));
    layer2_outputs(7961) <= layer1_outputs(8756);
    layer2_outputs(7962) <= not(layer1_outputs(10032)) or (layer1_outputs(7836));
    layer2_outputs(7963) <= (layer1_outputs(9362)) or (layer1_outputs(7871));
    layer2_outputs(7964) <= layer1_outputs(3825);
    layer2_outputs(7965) <= layer1_outputs(864);
    layer2_outputs(7966) <= layer1_outputs(4260);
    layer2_outputs(7967) <= (layer1_outputs(4995)) and not (layer1_outputs(4435));
    layer2_outputs(7968) <= not(layer1_outputs(3147)) or (layer1_outputs(9405));
    layer2_outputs(7969) <= not((layer1_outputs(2900)) or (layer1_outputs(7466)));
    layer2_outputs(7970) <= layer1_outputs(1216);
    layer2_outputs(7971) <= not(layer1_outputs(1910)) or (layer1_outputs(2256));
    layer2_outputs(7972) <= layer1_outputs(3912);
    layer2_outputs(7973) <= not(layer1_outputs(5472));
    layer2_outputs(7974) <= layer1_outputs(4384);
    layer2_outputs(7975) <= not(layer1_outputs(8242)) or (layer1_outputs(5189));
    layer2_outputs(7976) <= layer1_outputs(9244);
    layer2_outputs(7977) <= not(layer1_outputs(2440)) or (layer1_outputs(2676));
    layer2_outputs(7978) <= not((layer1_outputs(4726)) and (layer1_outputs(6553)));
    layer2_outputs(7979) <= not(layer1_outputs(6869));
    layer2_outputs(7980) <= layer1_outputs(2366);
    layer2_outputs(7981) <= not(layer1_outputs(10170));
    layer2_outputs(7982) <= layer1_outputs(4052);
    layer2_outputs(7983) <= layer1_outputs(956);
    layer2_outputs(7984) <= (layer1_outputs(8495)) or (layer1_outputs(8985));
    layer2_outputs(7985) <= '1';
    layer2_outputs(7986) <= layer1_outputs(8896);
    layer2_outputs(7987) <= (layer1_outputs(1112)) and not (layer1_outputs(7004));
    layer2_outputs(7988) <= (layer1_outputs(6381)) or (layer1_outputs(7914));
    layer2_outputs(7989) <= (layer1_outputs(8227)) and not (layer1_outputs(8213));
    layer2_outputs(7990) <= not((layer1_outputs(1642)) xor (layer1_outputs(5339)));
    layer2_outputs(7991) <= not((layer1_outputs(9794)) xor (layer1_outputs(7614)));
    layer2_outputs(7992) <= layer1_outputs(2117);
    layer2_outputs(7993) <= not(layer1_outputs(9609));
    layer2_outputs(7994) <= not(layer1_outputs(2859));
    layer2_outputs(7995) <= layer1_outputs(2449);
    layer2_outputs(7996) <= (layer1_outputs(6033)) and not (layer1_outputs(4127));
    layer2_outputs(7997) <= not((layer1_outputs(8305)) and (layer1_outputs(5047)));
    layer2_outputs(7998) <= (layer1_outputs(7660)) and not (layer1_outputs(1180));
    layer2_outputs(7999) <= not(layer1_outputs(9496));
    layer2_outputs(8000) <= (layer1_outputs(1534)) and (layer1_outputs(9641));
    layer2_outputs(8001) <= not(layer1_outputs(6452));
    layer2_outputs(8002) <= (layer1_outputs(6529)) xor (layer1_outputs(1566));
    layer2_outputs(8003) <= not(layer1_outputs(9537));
    layer2_outputs(8004) <= not(layer1_outputs(7907));
    layer2_outputs(8005) <= layer1_outputs(2138);
    layer2_outputs(8006) <= not((layer1_outputs(6164)) or (layer1_outputs(9957)));
    layer2_outputs(8007) <= (layer1_outputs(6934)) and not (layer1_outputs(5691));
    layer2_outputs(8008) <= not((layer1_outputs(731)) or (layer1_outputs(3993)));
    layer2_outputs(8009) <= (layer1_outputs(7182)) xor (layer1_outputs(3096));
    layer2_outputs(8010) <= layer1_outputs(3508);
    layer2_outputs(8011) <= (layer1_outputs(7106)) and not (layer1_outputs(578));
    layer2_outputs(8012) <= layer1_outputs(1729);
    layer2_outputs(8013) <= not(layer1_outputs(9566));
    layer2_outputs(8014) <= not(layer1_outputs(1146));
    layer2_outputs(8015) <= layer1_outputs(8466);
    layer2_outputs(8016) <= not((layer1_outputs(1771)) and (layer1_outputs(7953)));
    layer2_outputs(8017) <= (layer1_outputs(8589)) and not (layer1_outputs(4227));
    layer2_outputs(8018) <= (layer1_outputs(1178)) and not (layer1_outputs(1917));
    layer2_outputs(8019) <= (layer1_outputs(6317)) and not (layer1_outputs(1849));
    layer2_outputs(8020) <= (layer1_outputs(8113)) and not (layer1_outputs(1480));
    layer2_outputs(8021) <= not((layer1_outputs(6190)) and (layer1_outputs(6767)));
    layer2_outputs(8022) <= not((layer1_outputs(5727)) xor (layer1_outputs(6440)));
    layer2_outputs(8023) <= (layer1_outputs(6626)) xor (layer1_outputs(6720));
    layer2_outputs(8024) <= not((layer1_outputs(6210)) and (layer1_outputs(8474)));
    layer2_outputs(8025) <= (layer1_outputs(3483)) xor (layer1_outputs(10098));
    layer2_outputs(8026) <= not(layer1_outputs(4450));
    layer2_outputs(8027) <= not((layer1_outputs(6934)) or (layer1_outputs(1297)));
    layer2_outputs(8028) <= not(layer1_outputs(889));
    layer2_outputs(8029) <= not(layer1_outputs(3663));
    layer2_outputs(8030) <= (layer1_outputs(4546)) and not (layer1_outputs(492));
    layer2_outputs(8031) <= not(layer1_outputs(7552));
    layer2_outputs(8032) <= not((layer1_outputs(1771)) xor (layer1_outputs(7027)));
    layer2_outputs(8033) <= not(layer1_outputs(6376));
    layer2_outputs(8034) <= (layer1_outputs(4848)) and (layer1_outputs(7091));
    layer2_outputs(8035) <= not(layer1_outputs(8562)) or (layer1_outputs(3175));
    layer2_outputs(8036) <= (layer1_outputs(9672)) xor (layer1_outputs(9162));
    layer2_outputs(8037) <= layer1_outputs(2437);
    layer2_outputs(8038) <= layer1_outputs(2141);
    layer2_outputs(8039) <= not(layer1_outputs(756));
    layer2_outputs(8040) <= not(layer1_outputs(9339)) or (layer1_outputs(10058));
    layer2_outputs(8041) <= (layer1_outputs(5039)) xor (layer1_outputs(7097));
    layer2_outputs(8042) <= not(layer1_outputs(6400));
    layer2_outputs(8043) <= not(layer1_outputs(3722));
    layer2_outputs(8044) <= not(layer1_outputs(6559));
    layer2_outputs(8045) <= (layer1_outputs(2358)) or (layer1_outputs(5290));
    layer2_outputs(8046) <= not(layer1_outputs(8862)) or (layer1_outputs(9488));
    layer2_outputs(8047) <= layer1_outputs(124);
    layer2_outputs(8048) <= (layer1_outputs(1562)) and not (layer1_outputs(9968));
    layer2_outputs(8049) <= layer1_outputs(3507);
    layer2_outputs(8050) <= (layer1_outputs(1672)) and (layer1_outputs(3583));
    layer2_outputs(8051) <= layer1_outputs(9648);
    layer2_outputs(8052) <= not((layer1_outputs(7324)) or (layer1_outputs(2660)));
    layer2_outputs(8053) <= not(layer1_outputs(4578));
    layer2_outputs(8054) <= (layer1_outputs(7602)) and (layer1_outputs(4712));
    layer2_outputs(8055) <= (layer1_outputs(1265)) or (layer1_outputs(253));
    layer2_outputs(8056) <= not(layer1_outputs(6754));
    layer2_outputs(8057) <= not(layer1_outputs(4441));
    layer2_outputs(8058) <= (layer1_outputs(4792)) and not (layer1_outputs(9833));
    layer2_outputs(8059) <= (layer1_outputs(7242)) and not (layer1_outputs(2130));
    layer2_outputs(8060) <= (layer1_outputs(5024)) and not (layer1_outputs(3129));
    layer2_outputs(8061) <= not(layer1_outputs(9341));
    layer2_outputs(8062) <= not(layer1_outputs(349));
    layer2_outputs(8063) <= (layer1_outputs(7520)) or (layer1_outputs(3203));
    layer2_outputs(8064) <= not((layer1_outputs(2123)) or (layer1_outputs(9571)));
    layer2_outputs(8065) <= layer1_outputs(1418);
    layer2_outputs(8066) <= not(layer1_outputs(4619));
    layer2_outputs(8067) <= layer1_outputs(10183);
    layer2_outputs(8068) <= layer1_outputs(4154);
    layer2_outputs(8069) <= not((layer1_outputs(9687)) or (layer1_outputs(5009)));
    layer2_outputs(8070) <= not((layer1_outputs(8444)) and (layer1_outputs(6669)));
    layer2_outputs(8071) <= not((layer1_outputs(5832)) or (layer1_outputs(1318)));
    layer2_outputs(8072) <= layer1_outputs(2310);
    layer2_outputs(8073) <= (layer1_outputs(8839)) and (layer1_outputs(6299));
    layer2_outputs(8074) <= not(layer1_outputs(2140));
    layer2_outputs(8075) <= not(layer1_outputs(8929));
    layer2_outputs(8076) <= (layer1_outputs(809)) xor (layer1_outputs(6913));
    layer2_outputs(8077) <= not(layer1_outputs(4611));
    layer2_outputs(8078) <= not(layer1_outputs(5357));
    layer2_outputs(8079) <= not(layer1_outputs(2010));
    layer2_outputs(8080) <= not(layer1_outputs(4593));
    layer2_outputs(8081) <= not(layer1_outputs(1157));
    layer2_outputs(8082) <= not((layer1_outputs(8504)) and (layer1_outputs(9869)));
    layer2_outputs(8083) <= not(layer1_outputs(9213)) or (layer1_outputs(7466));
    layer2_outputs(8084) <= not(layer1_outputs(5767));
    layer2_outputs(8085) <= not(layer1_outputs(5815)) or (layer1_outputs(5626));
    layer2_outputs(8086) <= (layer1_outputs(8234)) xor (layer1_outputs(3638));
    layer2_outputs(8087) <= not((layer1_outputs(10218)) or (layer1_outputs(5616)));
    layer2_outputs(8088) <= not(layer1_outputs(8757));
    layer2_outputs(8089) <= not(layer1_outputs(6575));
    layer2_outputs(8090) <= not((layer1_outputs(4431)) and (layer1_outputs(3782)));
    layer2_outputs(8091) <= not(layer1_outputs(2086));
    layer2_outputs(8092) <= layer1_outputs(4629);
    layer2_outputs(8093) <= not(layer1_outputs(7832));
    layer2_outputs(8094) <= not(layer1_outputs(1082));
    layer2_outputs(8095) <= layer1_outputs(3883);
    layer2_outputs(8096) <= (layer1_outputs(6176)) and not (layer1_outputs(5418));
    layer2_outputs(8097) <= not(layer1_outputs(2913));
    layer2_outputs(8098) <= layer1_outputs(1974);
    layer2_outputs(8099) <= (layer1_outputs(8614)) or (layer1_outputs(3575));
    layer2_outputs(8100) <= (layer1_outputs(7450)) and not (layer1_outputs(4168));
    layer2_outputs(8101) <= layer1_outputs(4962);
    layer2_outputs(8102) <= not(layer1_outputs(10214));
    layer2_outputs(8103) <= not(layer1_outputs(3068)) or (layer1_outputs(6006));
    layer2_outputs(8104) <= not(layer1_outputs(9685));
    layer2_outputs(8105) <= not(layer1_outputs(6625));
    layer2_outputs(8106) <= not(layer1_outputs(8362));
    layer2_outputs(8107) <= (layer1_outputs(5258)) and not (layer1_outputs(9228));
    layer2_outputs(8108) <= layer1_outputs(10053);
    layer2_outputs(8109) <= (layer1_outputs(3532)) and not (layer1_outputs(2961));
    layer2_outputs(8110) <= (layer1_outputs(2587)) or (layer1_outputs(1092));
    layer2_outputs(8111) <= not(layer1_outputs(1219)) or (layer1_outputs(959));
    layer2_outputs(8112) <= (layer1_outputs(4040)) xor (layer1_outputs(6250));
    layer2_outputs(8113) <= not((layer1_outputs(797)) xor (layer1_outputs(7768)));
    layer2_outputs(8114) <= layer1_outputs(7788);
    layer2_outputs(8115) <= not(layer1_outputs(6507));
    layer2_outputs(8116) <= not(layer1_outputs(5932));
    layer2_outputs(8117) <= layer1_outputs(6965);
    layer2_outputs(8118) <= (layer1_outputs(10131)) xor (layer1_outputs(6154));
    layer2_outputs(8119) <= not(layer1_outputs(426));
    layer2_outputs(8120) <= not(layer1_outputs(3459));
    layer2_outputs(8121) <= (layer1_outputs(8963)) xor (layer1_outputs(2943));
    layer2_outputs(8122) <= not(layer1_outputs(9102));
    layer2_outputs(8123) <= (layer1_outputs(7483)) and not (layer1_outputs(2667));
    layer2_outputs(8124) <= not(layer1_outputs(7650));
    layer2_outputs(8125) <= (layer1_outputs(7714)) and not (layer1_outputs(620));
    layer2_outputs(8126) <= not(layer1_outputs(4221)) or (layer1_outputs(7174));
    layer2_outputs(8127) <= (layer1_outputs(9004)) xor (layer1_outputs(9590));
    layer2_outputs(8128) <= (layer1_outputs(3610)) and (layer1_outputs(1806));
    layer2_outputs(8129) <= (layer1_outputs(2397)) and (layer1_outputs(10237));
    layer2_outputs(8130) <= not(layer1_outputs(3539));
    layer2_outputs(8131) <= (layer1_outputs(9192)) and not (layer1_outputs(1475));
    layer2_outputs(8132) <= not(layer1_outputs(2946));
    layer2_outputs(8133) <= (layer1_outputs(9225)) or (layer1_outputs(7104));
    layer2_outputs(8134) <= (layer1_outputs(1818)) and (layer1_outputs(3277));
    layer2_outputs(8135) <= layer1_outputs(8133);
    layer2_outputs(8136) <= not(layer1_outputs(400));
    layer2_outputs(8137) <= not(layer1_outputs(5181));
    layer2_outputs(8138) <= not((layer1_outputs(3141)) and (layer1_outputs(6914)));
    layer2_outputs(8139) <= not(layer1_outputs(1671));
    layer2_outputs(8140) <= (layer1_outputs(8816)) and not (layer1_outputs(6829));
    layer2_outputs(8141) <= layer1_outputs(808);
    layer2_outputs(8142) <= not(layer1_outputs(8352)) or (layer1_outputs(1586));
    layer2_outputs(8143) <= not(layer1_outputs(5903)) or (layer1_outputs(6471));
    layer2_outputs(8144) <= layer1_outputs(3325);
    layer2_outputs(8145) <= (layer1_outputs(1535)) and not (layer1_outputs(9011));
    layer2_outputs(8146) <= not((layer1_outputs(4741)) or (layer1_outputs(4133)));
    layer2_outputs(8147) <= not((layer1_outputs(127)) xor (layer1_outputs(795)));
    layer2_outputs(8148) <= not(layer1_outputs(509)) or (layer1_outputs(5262));
    layer2_outputs(8149) <= layer1_outputs(236);
    layer2_outputs(8150) <= not(layer1_outputs(9673)) or (layer1_outputs(2246));
    layer2_outputs(8151) <= (layer1_outputs(4697)) and not (layer1_outputs(3436));
    layer2_outputs(8152) <= (layer1_outputs(7959)) or (layer1_outputs(7905));
    layer2_outputs(8153) <= (layer1_outputs(8354)) and not (layer1_outputs(6185));
    layer2_outputs(8154) <= (layer1_outputs(2460)) xor (layer1_outputs(8166));
    layer2_outputs(8155) <= not(layer1_outputs(1257));
    layer2_outputs(8156) <= (layer1_outputs(3688)) and (layer1_outputs(4124));
    layer2_outputs(8157) <= (layer1_outputs(372)) and (layer1_outputs(8544));
    layer2_outputs(8158) <= not((layer1_outputs(4601)) xor (layer1_outputs(1909)));
    layer2_outputs(8159) <= layer1_outputs(7717);
    layer2_outputs(8160) <= layer1_outputs(5054);
    layer2_outputs(8161) <= (layer1_outputs(161)) and (layer1_outputs(4905));
    layer2_outputs(8162) <= (layer1_outputs(8565)) and (layer1_outputs(4325));
    layer2_outputs(8163) <= not((layer1_outputs(3285)) or (layer1_outputs(3228)));
    layer2_outputs(8164) <= not(layer1_outputs(4941));
    layer2_outputs(8165) <= not(layer1_outputs(7589));
    layer2_outputs(8166) <= not(layer1_outputs(6473));
    layer2_outputs(8167) <= not(layer1_outputs(6595));
    layer2_outputs(8168) <= not(layer1_outputs(8571)) or (layer1_outputs(338));
    layer2_outputs(8169) <= (layer1_outputs(9674)) and not (layer1_outputs(5017));
    layer2_outputs(8170) <= not(layer1_outputs(3711));
    layer2_outputs(8171) <= (layer1_outputs(3142)) xor (layer1_outputs(5073));
    layer2_outputs(8172) <= not(layer1_outputs(1218));
    layer2_outputs(8173) <= not((layer1_outputs(6631)) and (layer1_outputs(6234)));
    layer2_outputs(8174) <= layer1_outputs(8465);
    layer2_outputs(8175) <= (layer1_outputs(7498)) and (layer1_outputs(4172));
    layer2_outputs(8176) <= layer1_outputs(5521);
    layer2_outputs(8177) <= (layer1_outputs(5146)) and not (layer1_outputs(4014));
    layer2_outputs(8178) <= not(layer1_outputs(3713));
    layer2_outputs(8179) <= (layer1_outputs(1557)) xor (layer1_outputs(7641));
    layer2_outputs(8180) <= not((layer1_outputs(1896)) and (layer1_outputs(4060)));
    layer2_outputs(8181) <= layer1_outputs(6546);
    layer2_outputs(8182) <= (layer1_outputs(6602)) xor (layer1_outputs(1547));
    layer2_outputs(8183) <= layer1_outputs(9309);
    layer2_outputs(8184) <= not(layer1_outputs(3015));
    layer2_outputs(8185) <= (layer1_outputs(5844)) xor (layer1_outputs(9049));
    layer2_outputs(8186) <= not(layer1_outputs(466));
    layer2_outputs(8187) <= not(layer1_outputs(2723));
    layer2_outputs(8188) <= not(layer1_outputs(1369));
    layer2_outputs(8189) <= (layer1_outputs(4371)) and not (layer1_outputs(1676));
    layer2_outputs(8190) <= not(layer1_outputs(3124));
    layer2_outputs(8191) <= layer1_outputs(1612);
    layer2_outputs(8192) <= (layer1_outputs(1841)) and not (layer1_outputs(7706));
    layer2_outputs(8193) <= not(layer1_outputs(7887));
    layer2_outputs(8194) <= not(layer1_outputs(7728));
    layer2_outputs(8195) <= (layer1_outputs(2661)) and not (layer1_outputs(2422));
    layer2_outputs(8196) <= layer1_outputs(4034);
    layer2_outputs(8197) <= not(layer1_outputs(9681)) or (layer1_outputs(9066));
    layer2_outputs(8198) <= not(layer1_outputs(7388));
    layer2_outputs(8199) <= layer1_outputs(2535);
    layer2_outputs(8200) <= not((layer1_outputs(304)) or (layer1_outputs(106)));
    layer2_outputs(8201) <= (layer1_outputs(7826)) xor (layer1_outputs(2204));
    layer2_outputs(8202) <= not(layer1_outputs(1881)) or (layer1_outputs(8810));
    layer2_outputs(8203) <= not((layer1_outputs(70)) xor (layer1_outputs(6767)));
    layer2_outputs(8204) <= layer1_outputs(1924);
    layer2_outputs(8205) <= (layer1_outputs(4967)) or (layer1_outputs(7277));
    layer2_outputs(8206) <= not(layer1_outputs(2948));
    layer2_outputs(8207) <= not(layer1_outputs(5751));
    layer2_outputs(8208) <= not(layer1_outputs(9053));
    layer2_outputs(8209) <= layer1_outputs(8615);
    layer2_outputs(8210) <= not(layer1_outputs(5863));
    layer2_outputs(8211) <= layer1_outputs(982);
    layer2_outputs(8212) <= not(layer1_outputs(1163));
    layer2_outputs(8213) <= layer1_outputs(5698);
    layer2_outputs(8214) <= not((layer1_outputs(3473)) or (layer1_outputs(8451)));
    layer2_outputs(8215) <= not(layer1_outputs(2498));
    layer2_outputs(8216) <= not(layer1_outputs(6254));
    layer2_outputs(8217) <= (layer1_outputs(8036)) xor (layer1_outputs(6707));
    layer2_outputs(8218) <= layer1_outputs(2415);
    layer2_outputs(8219) <= layer1_outputs(3948);
    layer2_outputs(8220) <= not((layer1_outputs(7930)) and (layer1_outputs(3667)));
    layer2_outputs(8221) <= layer1_outputs(7351);
    layer2_outputs(8222) <= not(layer1_outputs(2346));
    layer2_outputs(8223) <= layer1_outputs(690);
    layer2_outputs(8224) <= not(layer1_outputs(6136));
    layer2_outputs(8225) <= not(layer1_outputs(4762)) or (layer1_outputs(854));
    layer2_outputs(8226) <= not(layer1_outputs(3603));
    layer2_outputs(8227) <= (layer1_outputs(5297)) and not (layer1_outputs(9239));
    layer2_outputs(8228) <= not((layer1_outputs(2275)) and (layer1_outputs(5738)));
    layer2_outputs(8229) <= (layer1_outputs(6895)) and not (layer1_outputs(7037));
    layer2_outputs(8230) <= not(layer1_outputs(3718)) or (layer1_outputs(690));
    layer2_outputs(8231) <= layer1_outputs(8308);
    layer2_outputs(8232) <= not((layer1_outputs(9394)) or (layer1_outputs(10142)));
    layer2_outputs(8233) <= (layer1_outputs(3936)) or (layer1_outputs(7370));
    layer2_outputs(8234) <= layer1_outputs(1161);
    layer2_outputs(8235) <= layer1_outputs(4692);
    layer2_outputs(8236) <= (layer1_outputs(1806)) and not (layer1_outputs(5392));
    layer2_outputs(8237) <= layer1_outputs(1865);
    layer2_outputs(8238) <= layer1_outputs(728);
    layer2_outputs(8239) <= (layer1_outputs(3673)) or (layer1_outputs(6235));
    layer2_outputs(8240) <= layer1_outputs(8076);
    layer2_outputs(8241) <= layer1_outputs(176);
    layer2_outputs(8242) <= (layer1_outputs(8849)) xor (layer1_outputs(928));
    layer2_outputs(8243) <= not(layer1_outputs(1398));
    layer2_outputs(8244) <= (layer1_outputs(5494)) or (layer1_outputs(8861));
    layer2_outputs(8245) <= (layer1_outputs(4376)) or (layer1_outputs(4934));
    layer2_outputs(8246) <= (layer1_outputs(7824)) xor (layer1_outputs(8265));
    layer2_outputs(8247) <= (layer1_outputs(9725)) and (layer1_outputs(568));
    layer2_outputs(8248) <= (layer1_outputs(9216)) or (layer1_outputs(1938));
    layer2_outputs(8249) <= (layer1_outputs(5783)) and not (layer1_outputs(9651));
    layer2_outputs(8250) <= (layer1_outputs(2833)) or (layer1_outputs(6303));
    layer2_outputs(8251) <= layer1_outputs(6822);
    layer2_outputs(8252) <= layer1_outputs(8863);
    layer2_outputs(8253) <= (layer1_outputs(2877)) or (layer1_outputs(7309));
    layer2_outputs(8254) <= not(layer1_outputs(2038));
    layer2_outputs(8255) <= (layer1_outputs(8027)) and not (layer1_outputs(2156));
    layer2_outputs(8256) <= (layer1_outputs(1823)) and not (layer1_outputs(2924));
    layer2_outputs(8257) <= layer1_outputs(4849);
    layer2_outputs(8258) <= (layer1_outputs(7756)) or (layer1_outputs(4931));
    layer2_outputs(8259) <= not(layer1_outputs(1404));
    layer2_outputs(8260) <= not((layer1_outputs(3255)) xor (layer1_outputs(463)));
    layer2_outputs(8261) <= not(layer1_outputs(4583));
    layer2_outputs(8262) <= (layer1_outputs(5865)) xor (layer1_outputs(9194));
    layer2_outputs(8263) <= not(layer1_outputs(9077)) or (layer1_outputs(3877));
    layer2_outputs(8264) <= not(layer1_outputs(4231));
    layer2_outputs(8265) <= layer1_outputs(6569);
    layer2_outputs(8266) <= not(layer1_outputs(10163));
    layer2_outputs(8267) <= not(layer1_outputs(2614));
    layer2_outputs(8268) <= layer1_outputs(10059);
    layer2_outputs(8269) <= layer1_outputs(6437);
    layer2_outputs(8270) <= layer1_outputs(7325);
    layer2_outputs(8271) <= not((layer1_outputs(7658)) and (layer1_outputs(5689)));
    layer2_outputs(8272) <= not(layer1_outputs(4599));
    layer2_outputs(8273) <= (layer1_outputs(6806)) and not (layer1_outputs(7554));
    layer2_outputs(8274) <= layer1_outputs(7781);
    layer2_outputs(8275) <= not(layer1_outputs(5268));
    layer2_outputs(8276) <= not(layer1_outputs(6989));
    layer2_outputs(8277) <= layer1_outputs(5598);
    layer2_outputs(8278) <= layer1_outputs(4550);
    layer2_outputs(8279) <= not(layer1_outputs(2510));
    layer2_outputs(8280) <= not((layer1_outputs(5536)) and (layer1_outputs(8367)));
    layer2_outputs(8281) <= (layer1_outputs(1937)) or (layer1_outputs(4750));
    layer2_outputs(8282) <= (layer1_outputs(7108)) and not (layer1_outputs(1594));
    layer2_outputs(8283) <= layer1_outputs(8134);
    layer2_outputs(8284) <= (layer1_outputs(6920)) xor (layer1_outputs(605));
    layer2_outputs(8285) <= not((layer1_outputs(3242)) and (layer1_outputs(10236)));
    layer2_outputs(8286) <= not(layer1_outputs(444));
    layer2_outputs(8287) <= layer1_outputs(2133);
    layer2_outputs(8288) <= not(layer1_outputs(5070));
    layer2_outputs(8289) <= not(layer1_outputs(4051));
    layer2_outputs(8290) <= not((layer1_outputs(9318)) or (layer1_outputs(8198)));
    layer2_outputs(8291) <= layer1_outputs(9759);
    layer2_outputs(8292) <= (layer1_outputs(20)) or (layer1_outputs(7598));
    layer2_outputs(8293) <= layer1_outputs(2213);
    layer2_outputs(8294) <= (layer1_outputs(97)) xor (layer1_outputs(1328));
    layer2_outputs(8295) <= layer1_outputs(4409);
    layer2_outputs(8296) <= (layer1_outputs(2234)) xor (layer1_outputs(927));
    layer2_outputs(8297) <= layer1_outputs(8100);
    layer2_outputs(8298) <= not(layer1_outputs(5200));
    layer2_outputs(8299) <= not(layer1_outputs(2956));
    layer2_outputs(8300) <= layer1_outputs(1836);
    layer2_outputs(8301) <= not(layer1_outputs(8659));
    layer2_outputs(8302) <= layer1_outputs(5920);
    layer2_outputs(8303) <= layer1_outputs(7787);
    layer2_outputs(8304) <= not(layer1_outputs(8679));
    layer2_outputs(8305) <= (layer1_outputs(6968)) and not (layer1_outputs(7295));
    layer2_outputs(8306) <= layer1_outputs(4200);
    layer2_outputs(8307) <= layer1_outputs(10151);
    layer2_outputs(8308) <= not(layer1_outputs(6226));
    layer2_outputs(8309) <= layer1_outputs(7230);
    layer2_outputs(8310) <= not(layer1_outputs(8115));
    layer2_outputs(8311) <= (layer1_outputs(2138)) and (layer1_outputs(6501));
    layer2_outputs(8312) <= not(layer1_outputs(5196));
    layer2_outputs(8313) <= (layer1_outputs(746)) and not (layer1_outputs(1689));
    layer2_outputs(8314) <= layer1_outputs(4808);
    layer2_outputs(8315) <= not((layer1_outputs(8262)) xor (layer1_outputs(2183)));
    layer2_outputs(8316) <= not((layer1_outputs(7382)) xor (layer1_outputs(3409)));
    layer2_outputs(8317) <= not(layer1_outputs(1972)) or (layer1_outputs(2502));
    layer2_outputs(8318) <= not(layer1_outputs(1739));
    layer2_outputs(8319) <= layer1_outputs(1192);
    layer2_outputs(8320) <= layer1_outputs(4728);
    layer2_outputs(8321) <= not((layer1_outputs(2658)) and (layer1_outputs(9989)));
    layer2_outputs(8322) <= not(layer1_outputs(7624));
    layer2_outputs(8323) <= not(layer1_outputs(4135));
    layer2_outputs(8324) <= (layer1_outputs(3407)) or (layer1_outputs(5324));
    layer2_outputs(8325) <= not(layer1_outputs(4825)) or (layer1_outputs(8393));
    layer2_outputs(8326) <= not(layer1_outputs(8994)) or (layer1_outputs(1256));
    layer2_outputs(8327) <= layer1_outputs(4486);
    layer2_outputs(8328) <= layer1_outputs(7152);
    layer2_outputs(8329) <= not(layer1_outputs(5630)) or (layer1_outputs(4868));
    layer2_outputs(8330) <= (layer1_outputs(2706)) or (layer1_outputs(1943));
    layer2_outputs(8331) <= layer1_outputs(2129);
    layer2_outputs(8332) <= layer1_outputs(330);
    layer2_outputs(8333) <= (layer1_outputs(4321)) and not (layer1_outputs(991));
    layer2_outputs(8334) <= not(layer1_outputs(4294));
    layer2_outputs(8335) <= (layer1_outputs(2584)) and (layer1_outputs(4824));
    layer2_outputs(8336) <= (layer1_outputs(5574)) and not (layer1_outputs(1283));
    layer2_outputs(8337) <= not(layer1_outputs(152));
    layer2_outputs(8338) <= not(layer1_outputs(3377)) or (layer1_outputs(1330));
    layer2_outputs(8339) <= not((layer1_outputs(42)) xor (layer1_outputs(6565)));
    layer2_outputs(8340) <= (layer1_outputs(4053)) xor (layer1_outputs(7256));
    layer2_outputs(8341) <= layer1_outputs(7463);
    layer2_outputs(8342) <= not(layer1_outputs(6012));
    layer2_outputs(8343) <= not(layer1_outputs(3081));
    layer2_outputs(8344) <= not(layer1_outputs(2665)) or (layer1_outputs(1709));
    layer2_outputs(8345) <= not(layer1_outputs(4181));
    layer2_outputs(8346) <= (layer1_outputs(6588)) and not (layer1_outputs(916));
    layer2_outputs(8347) <= (layer1_outputs(4576)) and (layer1_outputs(6816));
    layer2_outputs(8348) <= not(layer1_outputs(9260));
    layer2_outputs(8349) <= not((layer1_outputs(8928)) or (layer1_outputs(6056)));
    layer2_outputs(8350) <= layer1_outputs(6898);
    layer2_outputs(8351) <= layer1_outputs(7514);
    layer2_outputs(8352) <= not((layer1_outputs(9257)) or (layer1_outputs(3661)));
    layer2_outputs(8353) <= (layer1_outputs(7452)) and (layer1_outputs(9230));
    layer2_outputs(8354) <= not(layer1_outputs(7873));
    layer2_outputs(8355) <= not(layer1_outputs(4205));
    layer2_outputs(8356) <= (layer1_outputs(1530)) and not (layer1_outputs(4468));
    layer2_outputs(8357) <= not(layer1_outputs(8691));
    layer2_outputs(8358) <= layer1_outputs(8880);
    layer2_outputs(8359) <= not((layer1_outputs(7088)) or (layer1_outputs(6443)));
    layer2_outputs(8360) <= not((layer1_outputs(8828)) xor (layer1_outputs(8101)));
    layer2_outputs(8361) <= (layer1_outputs(3095)) and not (layer1_outputs(9962));
    layer2_outputs(8362) <= not((layer1_outputs(9806)) and (layer1_outputs(1286)));
    layer2_outputs(8363) <= (layer1_outputs(585)) and not (layer1_outputs(9972));
    layer2_outputs(8364) <= not(layer1_outputs(3676));
    layer2_outputs(8365) <= not(layer1_outputs(6079));
    layer2_outputs(8366) <= (layer1_outputs(2857)) and not (layer1_outputs(6462));
    layer2_outputs(8367) <= (layer1_outputs(2403)) xor (layer1_outputs(1401));
    layer2_outputs(8368) <= (layer1_outputs(8186)) or (layer1_outputs(6271));
    layer2_outputs(8369) <= (layer1_outputs(550)) xor (layer1_outputs(10205));
    layer2_outputs(8370) <= (layer1_outputs(1671)) and not (layer1_outputs(4048));
    layer2_outputs(8371) <= layer1_outputs(1907);
    layer2_outputs(8372) <= (layer1_outputs(2850)) xor (layer1_outputs(6734));
    layer2_outputs(8373) <= (layer1_outputs(6368)) xor (layer1_outputs(2746));
    layer2_outputs(8374) <= layer1_outputs(4917);
    layer2_outputs(8375) <= not((layer1_outputs(7372)) xor (layer1_outputs(9690)));
    layer2_outputs(8376) <= (layer1_outputs(3521)) and not (layer1_outputs(5040));
    layer2_outputs(8377) <= (layer1_outputs(9698)) and (layer1_outputs(9054));
    layer2_outputs(8378) <= layer1_outputs(1700);
    layer2_outputs(8379) <= (layer1_outputs(8669)) and not (layer1_outputs(6084));
    layer2_outputs(8380) <= not(layer1_outputs(2486));
    layer2_outputs(8381) <= not(layer1_outputs(8768));
    layer2_outputs(8382) <= (layer1_outputs(1188)) and not (layer1_outputs(9304));
    layer2_outputs(8383) <= not(layer1_outputs(1828)) or (layer1_outputs(2795));
    layer2_outputs(8384) <= (layer1_outputs(4929)) and not (layer1_outputs(2730));
    layer2_outputs(8385) <= not(layer1_outputs(5550)) or (layer1_outputs(6619));
    layer2_outputs(8386) <= not(layer1_outputs(158));
    layer2_outputs(8387) <= (layer1_outputs(2652)) and not (layer1_outputs(2769));
    layer2_outputs(8388) <= (layer1_outputs(8680)) and (layer1_outputs(9924));
    layer2_outputs(8389) <= (layer1_outputs(2868)) and (layer1_outputs(2237));
    layer2_outputs(8390) <= not(layer1_outputs(5124));
    layer2_outputs(8391) <= not(layer1_outputs(7350)) or (layer1_outputs(10060));
    layer2_outputs(8392) <= (layer1_outputs(10191)) or (layer1_outputs(6900));
    layer2_outputs(8393) <= layer1_outputs(9115);
    layer2_outputs(8394) <= (layer1_outputs(4680)) xor (layer1_outputs(3395));
    layer2_outputs(8395) <= not(layer1_outputs(9177));
    layer2_outputs(8396) <= not(layer1_outputs(4871)) or (layer1_outputs(8008));
    layer2_outputs(8397) <= not(layer1_outputs(645));
    layer2_outputs(8398) <= layer1_outputs(6597);
    layer2_outputs(8399) <= layer1_outputs(7099);
    layer2_outputs(8400) <= not((layer1_outputs(4950)) or (layer1_outputs(10174)));
    layer2_outputs(8401) <= layer1_outputs(3972);
    layer2_outputs(8402) <= (layer1_outputs(2516)) and (layer1_outputs(6655));
    layer2_outputs(8403) <= (layer1_outputs(699)) and not (layer1_outputs(2914));
    layer2_outputs(8404) <= layer1_outputs(7531);
    layer2_outputs(8405) <= not((layer1_outputs(5355)) or (layer1_outputs(9026)));
    layer2_outputs(8406) <= (layer1_outputs(6855)) xor (layer1_outputs(2616));
    layer2_outputs(8407) <= not((layer1_outputs(5701)) or (layer1_outputs(2172)));
    layer2_outputs(8408) <= not((layer1_outputs(7090)) xor (layer1_outputs(5118)));
    layer2_outputs(8409) <= (layer1_outputs(9360)) and not (layer1_outputs(4460));
    layer2_outputs(8410) <= not((layer1_outputs(2390)) and (layer1_outputs(9175)));
    layer2_outputs(8411) <= not(layer1_outputs(5764));
    layer2_outputs(8412) <= not(layer1_outputs(8561));
    layer2_outputs(8413) <= layer1_outputs(9168);
    layer2_outputs(8414) <= (layer1_outputs(3729)) and not (layer1_outputs(7493));
    layer2_outputs(8415) <= not(layer1_outputs(1261));
    layer2_outputs(8416) <= (layer1_outputs(10146)) and not (layer1_outputs(7735));
    layer2_outputs(8417) <= not(layer1_outputs(6760)) or (layer1_outputs(3411));
    layer2_outputs(8418) <= layer1_outputs(8622);
    layer2_outputs(8419) <= (layer1_outputs(9038)) or (layer1_outputs(2737));
    layer2_outputs(8420) <= not(layer1_outputs(966));
    layer2_outputs(8421) <= (layer1_outputs(7193)) or (layer1_outputs(1345));
    layer2_outputs(8422) <= (layer1_outputs(573)) or (layer1_outputs(1801));
    layer2_outputs(8423) <= (layer1_outputs(5822)) or (layer1_outputs(8214));
    layer2_outputs(8424) <= not(layer1_outputs(4992)) or (layer1_outputs(6873));
    layer2_outputs(8425) <= not((layer1_outputs(10028)) and (layer1_outputs(9887)));
    layer2_outputs(8426) <= not((layer1_outputs(4509)) and (layer1_outputs(2743)));
    layer2_outputs(8427) <= not(layer1_outputs(948)) or (layer1_outputs(10110));
    layer2_outputs(8428) <= not((layer1_outputs(3887)) or (layer1_outputs(1402)));
    layer2_outputs(8429) <= not((layer1_outputs(6699)) and (layer1_outputs(8571)));
    layer2_outputs(8430) <= layer1_outputs(3923);
    layer2_outputs(8431) <= not((layer1_outputs(1186)) xor (layer1_outputs(2495)));
    layer2_outputs(8432) <= not((layer1_outputs(10047)) xor (layer1_outputs(3680)));
    layer2_outputs(8433) <= not(layer1_outputs(8314));
    layer2_outputs(8434) <= not((layer1_outputs(1897)) or (layer1_outputs(1429)));
    layer2_outputs(8435) <= not(layer1_outputs(1903));
    layer2_outputs(8436) <= not((layer1_outputs(5227)) and (layer1_outputs(1605)));
    layer2_outputs(8437) <= not(layer1_outputs(6593)) or (layer1_outputs(5063));
    layer2_outputs(8438) <= not(layer1_outputs(1531));
    layer2_outputs(8439) <= layer1_outputs(6249);
    layer2_outputs(8440) <= (layer1_outputs(1939)) or (layer1_outputs(8347));
    layer2_outputs(8441) <= not((layer1_outputs(8307)) and (layer1_outputs(8296)));
    layer2_outputs(8442) <= not(layer1_outputs(7474));
    layer2_outputs(8443) <= layer1_outputs(7174);
    layer2_outputs(8444) <= not(layer1_outputs(3418));
    layer2_outputs(8445) <= (layer1_outputs(545)) xor (layer1_outputs(489));
    layer2_outputs(8446) <= not(layer1_outputs(5905)) or (layer1_outputs(708));
    layer2_outputs(8447) <= layer1_outputs(3003);
    layer2_outputs(8448) <= not(layer1_outputs(2150)) or (layer1_outputs(6100));
    layer2_outputs(8449) <= layer1_outputs(773);
    layer2_outputs(8450) <= not((layer1_outputs(0)) xor (layer1_outputs(9015)));
    layer2_outputs(8451) <= not(layer1_outputs(4655));
    layer2_outputs(8452) <= not(layer1_outputs(119));
    layer2_outputs(8453) <= not((layer1_outputs(474)) xor (layer1_outputs(2113)));
    layer2_outputs(8454) <= layer1_outputs(9813);
    layer2_outputs(8455) <= (layer1_outputs(8579)) or (layer1_outputs(43));
    layer2_outputs(8456) <= not((layer1_outputs(447)) or (layer1_outputs(7155)));
    layer2_outputs(8457) <= (layer1_outputs(5220)) and (layer1_outputs(1905));
    layer2_outputs(8458) <= not(layer1_outputs(5732));
    layer2_outputs(8459) <= (layer1_outputs(8967)) or (layer1_outputs(3504));
    layer2_outputs(8460) <= not(layer1_outputs(3011)) or (layer1_outputs(2060));
    layer2_outputs(8461) <= not(layer1_outputs(6970));
    layer2_outputs(8462) <= '1';
    layer2_outputs(8463) <= (layer1_outputs(9917)) xor (layer1_outputs(6740));
    layer2_outputs(8464) <= not(layer1_outputs(6268));
    layer2_outputs(8465) <= layer1_outputs(2623);
    layer2_outputs(8466) <= (layer1_outputs(332)) xor (layer1_outputs(5904));
    layer2_outputs(8467) <= not(layer1_outputs(6359));
    layer2_outputs(8468) <= not((layer1_outputs(4547)) xor (layer1_outputs(7835)));
    layer2_outputs(8469) <= not((layer1_outputs(8560)) xor (layer1_outputs(647)));
    layer2_outputs(8470) <= not(layer1_outputs(545));
    layer2_outputs(8471) <= layer1_outputs(3769);
    layer2_outputs(8472) <= layer1_outputs(9551);
    layer2_outputs(8473) <= not(layer1_outputs(4012));
    layer2_outputs(8474) <= layer1_outputs(5494);
    layer2_outputs(8475) <= (layer1_outputs(3302)) xor (layer1_outputs(9096));
    layer2_outputs(8476) <= (layer1_outputs(4130)) and (layer1_outputs(4811));
    layer2_outputs(8477) <= not((layer1_outputs(8855)) and (layer1_outputs(9084)));
    layer2_outputs(8478) <= layer1_outputs(7856);
    layer2_outputs(8479) <= not((layer1_outputs(3777)) xor (layer1_outputs(1315)));
    layer2_outputs(8480) <= layer1_outputs(7442);
    layer2_outputs(8481) <= (layer1_outputs(877)) and not (layer1_outputs(8279));
    layer2_outputs(8482) <= not(layer1_outputs(6860)) or (layer1_outputs(2561));
    layer2_outputs(8483) <= not(layer1_outputs(4744));
    layer2_outputs(8484) <= layer1_outputs(7281);
    layer2_outputs(8485) <= not((layer1_outputs(9378)) xor (layer1_outputs(6602)));
    layer2_outputs(8486) <= not(layer1_outputs(356)) or (layer1_outputs(3115));
    layer2_outputs(8487) <= not((layer1_outputs(2303)) or (layer1_outputs(3939)));
    layer2_outputs(8488) <= not((layer1_outputs(9248)) xor (layer1_outputs(9857)));
    layer2_outputs(8489) <= not(layer1_outputs(5807)) or (layer1_outputs(2056));
    layer2_outputs(8490) <= not((layer1_outputs(5380)) and (layer1_outputs(1654)));
    layer2_outputs(8491) <= (layer1_outputs(867)) xor (layer1_outputs(6420));
    layer2_outputs(8492) <= not((layer1_outputs(6943)) or (layer1_outputs(8348)));
    layer2_outputs(8493) <= not(layer1_outputs(7192)) or (layer1_outputs(4802));
    layer2_outputs(8494) <= not(layer1_outputs(3957));
    layer2_outputs(8495) <= not(layer1_outputs(5428));
    layer2_outputs(8496) <= (layer1_outputs(2981)) xor (layer1_outputs(6510));
    layer2_outputs(8497) <= layer1_outputs(4877);
    layer2_outputs(8498) <= (layer1_outputs(7620)) and not (layer1_outputs(6415));
    layer2_outputs(8499) <= not(layer1_outputs(4609)) or (layer1_outputs(73));
    layer2_outputs(8500) <= layer1_outputs(7335);
    layer2_outputs(8501) <= (layer1_outputs(2651)) and not (layer1_outputs(8703));
    layer2_outputs(8502) <= not(layer1_outputs(447));
    layer2_outputs(8503) <= (layer1_outputs(2049)) and not (layer1_outputs(2384));
    layer2_outputs(8504) <= not((layer1_outputs(3088)) xor (layer1_outputs(917)));
    layer2_outputs(8505) <= not(layer1_outputs(8705));
    layer2_outputs(8506) <= '0';
    layer2_outputs(8507) <= not(layer1_outputs(8637));
    layer2_outputs(8508) <= (layer1_outputs(467)) and (layer1_outputs(4492));
    layer2_outputs(8509) <= not((layer1_outputs(8352)) and (layer1_outputs(1941)));
    layer2_outputs(8510) <= (layer1_outputs(4829)) and not (layer1_outputs(6267));
    layer2_outputs(8511) <= not(layer1_outputs(4649));
    layer2_outputs(8512) <= not((layer1_outputs(2246)) and (layer1_outputs(8435)));
    layer2_outputs(8513) <= not(layer1_outputs(9397));
    layer2_outputs(8514) <= not(layer1_outputs(9090)) or (layer1_outputs(3025));
    layer2_outputs(8515) <= layer1_outputs(138);
    layer2_outputs(8516) <= layer1_outputs(7219);
    layer2_outputs(8517) <= (layer1_outputs(2387)) and not (layer1_outputs(474));
    layer2_outputs(8518) <= not((layer1_outputs(3622)) or (layer1_outputs(2513)));
    layer2_outputs(8519) <= layer1_outputs(7643);
    layer2_outputs(8520) <= (layer1_outputs(9161)) and not (layer1_outputs(409));
    layer2_outputs(8521) <= layer1_outputs(4350);
    layer2_outputs(8522) <= not((layer1_outputs(6555)) or (layer1_outputs(7467)));
    layer2_outputs(8523) <= layer1_outputs(8478);
    layer2_outputs(8524) <= not(layer1_outputs(630)) or (layer1_outputs(4304));
    layer2_outputs(8525) <= not((layer1_outputs(3175)) or (layer1_outputs(7742)));
    layer2_outputs(8526) <= layer1_outputs(3546);
    layer2_outputs(8527) <= not(layer1_outputs(9469));
    layer2_outputs(8528) <= not(layer1_outputs(2222));
    layer2_outputs(8529) <= (layer1_outputs(2848)) or (layer1_outputs(8311));
    layer2_outputs(8530) <= not(layer1_outputs(9312));
    layer2_outputs(8531) <= layer1_outputs(5252);
    layer2_outputs(8532) <= not((layer1_outputs(8941)) xor (layer1_outputs(7832)));
    layer2_outputs(8533) <= not(layer1_outputs(1316));
    layer2_outputs(8534) <= not((layer1_outputs(7547)) or (layer1_outputs(7181)));
    layer2_outputs(8535) <= not(layer1_outputs(311));
    layer2_outputs(8536) <= not(layer1_outputs(390));
    layer2_outputs(8537) <= not(layer1_outputs(3726));
    layer2_outputs(8538) <= (layer1_outputs(7344)) and (layer1_outputs(224));
    layer2_outputs(8539) <= layer1_outputs(8587);
    layer2_outputs(8540) <= not(layer1_outputs(1172));
    layer2_outputs(8541) <= not((layer1_outputs(674)) xor (layer1_outputs(8949)));
    layer2_outputs(8542) <= (layer1_outputs(5099)) or (layer1_outputs(3293));
    layer2_outputs(8543) <= layer1_outputs(1303);
    layer2_outputs(8544) <= '0';
    layer2_outputs(8545) <= layer1_outputs(3176);
    layer2_outputs(8546) <= not((layer1_outputs(7331)) or (layer1_outputs(9365)));
    layer2_outputs(8547) <= (layer1_outputs(6019)) or (layer1_outputs(5671));
    layer2_outputs(8548) <= not(layer1_outputs(2348)) or (layer1_outputs(9578));
    layer2_outputs(8549) <= layer1_outputs(5918);
    layer2_outputs(8550) <= not(layer1_outputs(1716));
    layer2_outputs(8551) <= (layer1_outputs(3647)) and (layer1_outputs(992));
    layer2_outputs(8552) <= (layer1_outputs(10)) or (layer1_outputs(3097));
    layer2_outputs(8553) <= (layer1_outputs(4259)) and not (layer1_outputs(7303));
    layer2_outputs(8554) <= not(layer1_outputs(1230));
    layer2_outputs(8555) <= not((layer1_outputs(8114)) and (layer1_outputs(2896)));
    layer2_outputs(8556) <= not(layer1_outputs(5187));
    layer2_outputs(8557) <= (layer1_outputs(3305)) and (layer1_outputs(5910));
    layer2_outputs(8558) <= not((layer1_outputs(1331)) xor (layer1_outputs(4259)));
    layer2_outputs(8559) <= not(layer1_outputs(80));
    layer2_outputs(8560) <= not(layer1_outputs(5537));
    layer2_outputs(8561) <= (layer1_outputs(1043)) xor (layer1_outputs(6001));
    layer2_outputs(8562) <= (layer1_outputs(8316)) and not (layer1_outputs(1329));
    layer2_outputs(8563) <= not(layer1_outputs(8428));
    layer2_outputs(8564) <= not(layer1_outputs(3044));
    layer2_outputs(8565) <= not(layer1_outputs(3108));
    layer2_outputs(8566) <= not(layer1_outputs(4709)) or (layer1_outputs(4757));
    layer2_outputs(8567) <= not(layer1_outputs(1528));
    layer2_outputs(8568) <= (layer1_outputs(7405)) and not (layer1_outputs(7846));
    layer2_outputs(8569) <= layer1_outputs(2944);
    layer2_outputs(8570) <= not(layer1_outputs(2477)) or (layer1_outputs(208));
    layer2_outputs(8571) <= (layer1_outputs(5700)) and not (layer1_outputs(9215));
    layer2_outputs(8572) <= layer1_outputs(6664);
    layer2_outputs(8573) <= not((layer1_outputs(5018)) or (layer1_outputs(2499)));
    layer2_outputs(8574) <= not((layer1_outputs(6646)) xor (layer1_outputs(2088)));
    layer2_outputs(8575) <= (layer1_outputs(9253)) and not (layer1_outputs(1287));
    layer2_outputs(8576) <= (layer1_outputs(595)) or (layer1_outputs(9965));
    layer2_outputs(8577) <= layer1_outputs(1128);
    layer2_outputs(8578) <= not(layer1_outputs(2051)) or (layer1_outputs(2101));
    layer2_outputs(8579) <= (layer1_outputs(9836)) or (layer1_outputs(1215));
    layer2_outputs(8580) <= (layer1_outputs(6983)) or (layer1_outputs(5703));
    layer2_outputs(8581) <= not(layer1_outputs(7374));
    layer2_outputs(8582) <= not(layer1_outputs(6043));
    layer2_outputs(8583) <= not(layer1_outputs(3052)) or (layer1_outputs(7253));
    layer2_outputs(8584) <= not(layer1_outputs(8925));
    layer2_outputs(8585) <= not(layer1_outputs(7285));
    layer2_outputs(8586) <= not(layer1_outputs(8724));
    layer2_outputs(8587) <= not(layer1_outputs(9914)) or (layer1_outputs(8959));
    layer2_outputs(8588) <= not(layer1_outputs(3953));
    layer2_outputs(8589) <= not(layer1_outputs(5560));
    layer2_outputs(8590) <= not(layer1_outputs(9110)) or (layer1_outputs(7982));
    layer2_outputs(8591) <= not(layer1_outputs(6508));
    layer2_outputs(8592) <= layer1_outputs(10109);
    layer2_outputs(8593) <= layer1_outputs(282);
    layer2_outputs(8594) <= not(layer1_outputs(6854));
    layer2_outputs(8595) <= (layer1_outputs(9377)) or (layer1_outputs(6404));
    layer2_outputs(8596) <= not(layer1_outputs(1600));
    layer2_outputs(8597) <= not((layer1_outputs(5469)) and (layer1_outputs(9136)));
    layer2_outputs(8598) <= (layer1_outputs(5712)) xor (layer1_outputs(773));
    layer2_outputs(8599) <= not(layer1_outputs(7109)) or (layer1_outputs(2531));
    layer2_outputs(8600) <= not((layer1_outputs(9669)) and (layer1_outputs(2629)));
    layer2_outputs(8601) <= (layer1_outputs(9279)) xor (layer1_outputs(7570));
    layer2_outputs(8602) <= not(layer1_outputs(3605));
    layer2_outputs(8603) <= (layer1_outputs(9921)) xor (layer1_outputs(847));
    layer2_outputs(8604) <= not(layer1_outputs(9677)) or (layer1_outputs(5985));
    layer2_outputs(8605) <= layer1_outputs(6844);
    layer2_outputs(8606) <= not(layer1_outputs(7502)) or (layer1_outputs(677));
    layer2_outputs(8607) <= (layer1_outputs(4169)) or (layer1_outputs(7897));
    layer2_outputs(8608) <= layer1_outputs(9024);
    layer2_outputs(8609) <= (layer1_outputs(6857)) and (layer1_outputs(7901));
    layer2_outputs(8610) <= not(layer1_outputs(1784));
    layer2_outputs(8611) <= not(layer1_outputs(8475));
    layer2_outputs(8612) <= not(layer1_outputs(1046));
    layer2_outputs(8613) <= not(layer1_outputs(6486));
    layer2_outputs(8614) <= (layer1_outputs(2697)) and (layer1_outputs(1053));
    layer2_outputs(8615) <= layer1_outputs(6889);
    layer2_outputs(8616) <= layer1_outputs(9280);
    layer2_outputs(8617) <= layer1_outputs(5718);
    layer2_outputs(8618) <= (layer1_outputs(351)) and (layer1_outputs(1708));
    layer2_outputs(8619) <= (layer1_outputs(2121)) and (layer1_outputs(5635));
    layer2_outputs(8620) <= not((layer1_outputs(8072)) or (layer1_outputs(6994)));
    layer2_outputs(8621) <= not(layer1_outputs(3788));
    layer2_outputs(8622) <= not(layer1_outputs(126)) or (layer1_outputs(8981));
    layer2_outputs(8623) <= not((layer1_outputs(744)) or (layer1_outputs(9471)));
    layer2_outputs(8624) <= layer1_outputs(5453);
    layer2_outputs(8625) <= not(layer1_outputs(2170));
    layer2_outputs(8626) <= not(layer1_outputs(2087));
    layer2_outputs(8627) <= (layer1_outputs(5759)) or (layer1_outputs(4374));
    layer2_outputs(8628) <= layer1_outputs(3352);
    layer2_outputs(8629) <= (layer1_outputs(7536)) and not (layer1_outputs(8361));
    layer2_outputs(8630) <= layer1_outputs(8092);
    layer2_outputs(8631) <= (layer1_outputs(2757)) or (layer1_outputs(46));
    layer2_outputs(8632) <= not((layer1_outputs(7879)) xor (layer1_outputs(6450)));
    layer2_outputs(8633) <= not((layer1_outputs(4870)) and (layer1_outputs(9657)));
    layer2_outputs(8634) <= (layer1_outputs(5948)) xor (layer1_outputs(6769));
    layer2_outputs(8635) <= (layer1_outputs(7394)) or (layer1_outputs(44));
    layer2_outputs(8636) <= not(layer1_outputs(242)) or (layer1_outputs(8115));
    layer2_outputs(8637) <= not(layer1_outputs(4460));
    layer2_outputs(8638) <= '1';
    layer2_outputs(8639) <= not((layer1_outputs(7854)) xor (layer1_outputs(2625)));
    layer2_outputs(8640) <= (layer1_outputs(8644)) xor (layer1_outputs(3673));
    layer2_outputs(8641) <= not(layer1_outputs(1610)) or (layer1_outputs(5140));
    layer2_outputs(8642) <= not((layer1_outputs(4287)) xor (layer1_outputs(4747)));
    layer2_outputs(8643) <= layer1_outputs(5594);
    layer2_outputs(8644) <= (layer1_outputs(8673)) xor (layer1_outputs(844));
    layer2_outputs(8645) <= not((layer1_outputs(4278)) and (layer1_outputs(4552)));
    layer2_outputs(8646) <= not((layer1_outputs(5312)) and (layer1_outputs(3487)));
    layer2_outputs(8647) <= not((layer1_outputs(4935)) and (layer1_outputs(5951)));
    layer2_outputs(8648) <= (layer1_outputs(4816)) and not (layer1_outputs(8872));
    layer2_outputs(8649) <= not(layer1_outputs(3000));
    layer2_outputs(8650) <= (layer1_outputs(6207)) and (layer1_outputs(3712));
    layer2_outputs(8651) <= not(layer1_outputs(7902));
    layer2_outputs(8652) <= (layer1_outputs(2897)) xor (layer1_outputs(8326));
    layer2_outputs(8653) <= not(layer1_outputs(6085));
    layer2_outputs(8654) <= not((layer1_outputs(5557)) and (layer1_outputs(7537)));
    layer2_outputs(8655) <= '1';
    layer2_outputs(8656) <= not(layer1_outputs(6302));
    layer2_outputs(8657) <= (layer1_outputs(2563)) and not (layer1_outputs(9358));
    layer2_outputs(8658) <= layer1_outputs(8019);
    layer2_outputs(8659) <= not(layer1_outputs(9544)) or (layer1_outputs(6568));
    layer2_outputs(8660) <= layer1_outputs(10056);
    layer2_outputs(8661) <= not((layer1_outputs(9297)) and (layer1_outputs(6560)));
    layer2_outputs(8662) <= layer1_outputs(133);
    layer2_outputs(8663) <= not(layer1_outputs(6650));
    layer2_outputs(8664) <= (layer1_outputs(5126)) xor (layer1_outputs(8785));
    layer2_outputs(8665) <= not((layer1_outputs(4267)) and (layer1_outputs(3771)));
    layer2_outputs(8666) <= layer1_outputs(4862);
    layer2_outputs(8667) <= not(layer1_outputs(3813));
    layer2_outputs(8668) <= not((layer1_outputs(1734)) and (layer1_outputs(5132)));
    layer2_outputs(8669) <= not(layer1_outputs(884));
    layer2_outputs(8670) <= (layer1_outputs(7298)) xor (layer1_outputs(9927));
    layer2_outputs(8671) <= not(layer1_outputs(2926));
    layer2_outputs(8672) <= (layer1_outputs(3346)) xor (layer1_outputs(3364));
    layer2_outputs(8673) <= layer1_outputs(6386);
    layer2_outputs(8674) <= (layer1_outputs(4809)) xor (layer1_outputs(8764));
    layer2_outputs(8675) <= not(layer1_outputs(6736));
    layer2_outputs(8676) <= layer1_outputs(7727);
    layer2_outputs(8677) <= (layer1_outputs(624)) or (layer1_outputs(2333));
    layer2_outputs(8678) <= layer1_outputs(518);
    layer2_outputs(8679) <= layer1_outputs(7899);
    layer2_outputs(8680) <= '1';
    layer2_outputs(8681) <= layer1_outputs(10211);
    layer2_outputs(8682) <= not(layer1_outputs(3840));
    layer2_outputs(8683) <= layer1_outputs(4109);
    layer2_outputs(8684) <= (layer1_outputs(4617)) or (layer1_outputs(3720));
    layer2_outputs(8685) <= (layer1_outputs(6708)) and not (layer1_outputs(1452));
    layer2_outputs(8686) <= layer1_outputs(5188);
    layer2_outputs(8687) <= not(layer1_outputs(10003));
    layer2_outputs(8688) <= (layer1_outputs(8637)) or (layer1_outputs(6909));
    layer2_outputs(8689) <= not(layer1_outputs(4254));
    layer2_outputs(8690) <= (layer1_outputs(2128)) and not (layer1_outputs(1098));
    layer2_outputs(8691) <= not(layer1_outputs(9211));
    layer2_outputs(8692) <= layer1_outputs(315);
    layer2_outputs(8693) <= '0';
    layer2_outputs(8694) <= (layer1_outputs(3389)) and not (layer1_outputs(3341));
    layer2_outputs(8695) <= layer1_outputs(10113);
    layer2_outputs(8696) <= not(layer1_outputs(93));
    layer2_outputs(8697) <= (layer1_outputs(8790)) xor (layer1_outputs(3391));
    layer2_outputs(8698) <= not((layer1_outputs(4968)) xor (layer1_outputs(5928)));
    layer2_outputs(8699) <= layer1_outputs(3969);
    layer2_outputs(8700) <= not(layer1_outputs(1961)) or (layer1_outputs(176));
    layer2_outputs(8701) <= not((layer1_outputs(6864)) or (layer1_outputs(3770)));
    layer2_outputs(8702) <= layer1_outputs(10223);
    layer2_outputs(8703) <= layer1_outputs(1015);
    layer2_outputs(8704) <= not(layer1_outputs(3472)) or (layer1_outputs(9030));
    layer2_outputs(8705) <= not(layer1_outputs(7950));
    layer2_outputs(8706) <= layer1_outputs(3589);
    layer2_outputs(8707) <= layer1_outputs(3286);
    layer2_outputs(8708) <= layer1_outputs(238);
    layer2_outputs(8709) <= not(layer1_outputs(8044));
    layer2_outputs(8710) <= (layer1_outputs(7787)) xor (layer1_outputs(10193));
    layer2_outputs(8711) <= (layer1_outputs(8088)) and not (layer1_outputs(8397));
    layer2_outputs(8712) <= not(layer1_outputs(9741));
    layer2_outputs(8713) <= not(layer1_outputs(9848));
    layer2_outputs(8714) <= not(layer1_outputs(273));
    layer2_outputs(8715) <= not(layer1_outputs(4801));
    layer2_outputs(8716) <= (layer1_outputs(25)) or (layer1_outputs(1481));
    layer2_outputs(8717) <= (layer1_outputs(9623)) and not (layer1_outputs(6451));
    layer2_outputs(8718) <= not(layer1_outputs(3368));
    layer2_outputs(8719) <= not(layer1_outputs(5069));
    layer2_outputs(8720) <= not((layer1_outputs(9877)) and (layer1_outputs(1790)));
    layer2_outputs(8721) <= not(layer1_outputs(10134));
    layer2_outputs(8722) <= layer1_outputs(9294);
    layer2_outputs(8723) <= (layer1_outputs(3794)) xor (layer1_outputs(1755));
    layer2_outputs(8724) <= layer1_outputs(8726);
    layer2_outputs(8725) <= (layer1_outputs(9730)) and (layer1_outputs(1570));
    layer2_outputs(8726) <= (layer1_outputs(8727)) and (layer1_outputs(8237));
    layer2_outputs(8727) <= layer1_outputs(532);
    layer2_outputs(8728) <= not(layer1_outputs(8013)) or (layer1_outputs(8740));
    layer2_outputs(8729) <= layer1_outputs(7609);
    layer2_outputs(8730) <= not(layer1_outputs(20));
    layer2_outputs(8731) <= not(layer1_outputs(6020)) or (layer1_outputs(7528));
    layer2_outputs(8732) <= layer1_outputs(3028);
    layer2_outputs(8733) <= layer1_outputs(10133);
    layer2_outputs(8734) <= layer1_outputs(5138);
    layer2_outputs(8735) <= not(layer1_outputs(637));
    layer2_outputs(8736) <= layer1_outputs(7270);
    layer2_outputs(8737) <= not(layer1_outputs(189));
    layer2_outputs(8738) <= layer1_outputs(8208);
    layer2_outputs(8739) <= (layer1_outputs(892)) or (layer1_outputs(6831));
    layer2_outputs(8740) <= layer1_outputs(905);
    layer2_outputs(8741) <= layer1_outputs(9529);
    layer2_outputs(8742) <= (layer1_outputs(10092)) and not (layer1_outputs(3449));
    layer2_outputs(8743) <= layer1_outputs(3949);
    layer2_outputs(8744) <= layer1_outputs(9151);
    layer2_outputs(8745) <= layer1_outputs(6189);
    layer2_outputs(8746) <= layer1_outputs(4197);
    layer2_outputs(8747) <= not(layer1_outputs(6980));
    layer2_outputs(8748) <= layer1_outputs(3131);
    layer2_outputs(8749) <= layer1_outputs(10231);
    layer2_outputs(8750) <= layer1_outputs(3979);
    layer2_outputs(8751) <= (layer1_outputs(6283)) and (layer1_outputs(4276));
    layer2_outputs(8752) <= (layer1_outputs(8849)) and not (layer1_outputs(3000));
    layer2_outputs(8753) <= not((layer1_outputs(3351)) or (layer1_outputs(9455)));
    layer2_outputs(8754) <= layer1_outputs(5301);
    layer2_outputs(8755) <= not(layer1_outputs(5007)) or (layer1_outputs(3946));
    layer2_outputs(8756) <= (layer1_outputs(6906)) and not (layer1_outputs(2565));
    layer2_outputs(8757) <= not(layer1_outputs(9067));
    layer2_outputs(8758) <= layer1_outputs(8798);
    layer2_outputs(8759) <= layer1_outputs(2990);
    layer2_outputs(8760) <= not(layer1_outputs(4688));
    layer2_outputs(8761) <= layer1_outputs(9509);
    layer2_outputs(8762) <= not(layer1_outputs(6118)) or (layer1_outputs(1745));
    layer2_outputs(8763) <= (layer1_outputs(3938)) and not (layer1_outputs(8089));
    layer2_outputs(8764) <= layer1_outputs(8908);
    layer2_outputs(8765) <= not(layer1_outputs(5184));
    layer2_outputs(8766) <= layer1_outputs(6471);
    layer2_outputs(8767) <= not((layer1_outputs(9767)) and (layer1_outputs(5138)));
    layer2_outputs(8768) <= layer1_outputs(10198);
    layer2_outputs(8769) <= not((layer1_outputs(7562)) xor (layer1_outputs(9033)));
    layer2_outputs(8770) <= not((layer1_outputs(3468)) xor (layer1_outputs(35)));
    layer2_outputs(8771) <= not(layer1_outputs(9234));
    layer2_outputs(8772) <= not(layer1_outputs(738));
    layer2_outputs(8773) <= layer1_outputs(464);
    layer2_outputs(8774) <= layer1_outputs(9567);
    layer2_outputs(8775) <= layer1_outputs(7028);
    layer2_outputs(8776) <= layer1_outputs(7230);
    layer2_outputs(8777) <= layer1_outputs(6264);
    layer2_outputs(8778) <= layer1_outputs(273);
    layer2_outputs(8779) <= not(layer1_outputs(1292)) or (layer1_outputs(1173));
    layer2_outputs(8780) <= not(layer1_outputs(8688));
    layer2_outputs(8781) <= layer1_outputs(2934);
    layer2_outputs(8782) <= not(layer1_outputs(5459));
    layer2_outputs(8783) <= not(layer1_outputs(946));
    layer2_outputs(8784) <= layer1_outputs(9916);
    layer2_outputs(8785) <= layer1_outputs(4036);
    layer2_outputs(8786) <= layer1_outputs(7546);
    layer2_outputs(8787) <= not(layer1_outputs(8558)) or (layer1_outputs(7562));
    layer2_outputs(8788) <= not(layer1_outputs(3711));
    layer2_outputs(8789) <= not((layer1_outputs(231)) xor (layer1_outputs(6124)));
    layer2_outputs(8790) <= not(layer1_outputs(8422));
    layer2_outputs(8791) <= not((layer1_outputs(6097)) and (layer1_outputs(4816)));
    layer2_outputs(8792) <= not(layer1_outputs(2366));
    layer2_outputs(8793) <= not(layer1_outputs(4894));
    layer2_outputs(8794) <= layer1_outputs(4865);
    layer2_outputs(8795) <= layer1_outputs(9068);
    layer2_outputs(8796) <= not(layer1_outputs(1495));
    layer2_outputs(8797) <= layer1_outputs(4517);
    layer2_outputs(8798) <= not(layer1_outputs(66));
    layer2_outputs(8799) <= (layer1_outputs(9850)) xor (layer1_outputs(6896));
    layer2_outputs(8800) <= not((layer1_outputs(4793)) xor (layer1_outputs(356)));
    layer2_outputs(8801) <= not(layer1_outputs(6198));
    layer2_outputs(8802) <= not((layer1_outputs(5605)) xor (layer1_outputs(3153)));
    layer2_outputs(8803) <= layer1_outputs(9270);
    layer2_outputs(8804) <= not((layer1_outputs(6237)) and (layer1_outputs(9754)));
    layer2_outputs(8805) <= not((layer1_outputs(3425)) and (layer1_outputs(1504)));
    layer2_outputs(8806) <= (layer1_outputs(7973)) xor (layer1_outputs(8586));
    layer2_outputs(8807) <= layer1_outputs(4684);
    layer2_outputs(8808) <= not(layer1_outputs(8038));
    layer2_outputs(8809) <= (layer1_outputs(3220)) or (layer1_outputs(8407));
    layer2_outputs(8810) <= (layer1_outputs(7188)) or (layer1_outputs(9902));
    layer2_outputs(8811) <= (layer1_outputs(1414)) or (layer1_outputs(9575));
    layer2_outputs(8812) <= not(layer1_outputs(4465));
    layer2_outputs(8813) <= not((layer1_outputs(856)) xor (layer1_outputs(3159)));
    layer2_outputs(8814) <= not((layer1_outputs(2719)) xor (layer1_outputs(2888)));
    layer2_outputs(8815) <= not(layer1_outputs(3577)) or (layer1_outputs(2910));
    layer2_outputs(8816) <= not(layer1_outputs(5345)) or (layer1_outputs(4521));
    layer2_outputs(8817) <= (layer1_outputs(10108)) and not (layer1_outputs(7640));
    layer2_outputs(8818) <= (layer1_outputs(8460)) and (layer1_outputs(5508));
    layer2_outputs(8819) <= not(layer1_outputs(6644));
    layer2_outputs(8820) <= not((layer1_outputs(4707)) xor (layer1_outputs(232)));
    layer2_outputs(8821) <= not(layer1_outputs(7178));
    layer2_outputs(8822) <= not((layer1_outputs(9692)) or (layer1_outputs(5327)));
    layer2_outputs(8823) <= (layer1_outputs(5275)) and not (layer1_outputs(2151));
    layer2_outputs(8824) <= layer1_outputs(7103);
    layer2_outputs(8825) <= not(layer1_outputs(3420));
    layer2_outputs(8826) <= (layer1_outputs(755)) and not (layer1_outputs(1945));
    layer2_outputs(8827) <= not((layer1_outputs(4957)) and (layer1_outputs(10194)));
    layer2_outputs(8828) <= not(layer1_outputs(5657)) or (layer1_outputs(4041));
    layer2_outputs(8829) <= layer1_outputs(6739);
    layer2_outputs(8830) <= layer1_outputs(2481);
    layer2_outputs(8831) <= (layer1_outputs(2956)) and not (layer1_outputs(2221));
    layer2_outputs(8832) <= layer1_outputs(335);
    layer2_outputs(8833) <= layer1_outputs(1911);
    layer2_outputs(8834) <= (layer1_outputs(4033)) and not (layer1_outputs(5434));
    layer2_outputs(8835) <= (layer1_outputs(5201)) and (layer1_outputs(4372));
    layer2_outputs(8836) <= not(layer1_outputs(824));
    layer2_outputs(8837) <= not((layer1_outputs(4558)) and (layer1_outputs(8907)));
    layer2_outputs(8838) <= (layer1_outputs(2083)) and not (layer1_outputs(4597));
    layer2_outputs(8839) <= not(layer1_outputs(5015));
    layer2_outputs(8840) <= not(layer1_outputs(7702));
    layer2_outputs(8841) <= (layer1_outputs(7432)) and not (layer1_outputs(8463));
    layer2_outputs(8842) <= not(layer1_outputs(1497));
    layer2_outputs(8843) <= not((layer1_outputs(1247)) or (layer1_outputs(8491)));
    layer2_outputs(8844) <= layer1_outputs(4640);
    layer2_outputs(8845) <= layer1_outputs(3990);
    layer2_outputs(8846) <= not(layer1_outputs(5655)) or (layer1_outputs(2585));
    layer2_outputs(8847) <= not(layer1_outputs(4592));
    layer2_outputs(8848) <= not(layer1_outputs(5819));
    layer2_outputs(8849) <= not(layer1_outputs(8010));
    layer2_outputs(8850) <= not(layer1_outputs(9574));
    layer2_outputs(8851) <= (layer1_outputs(6954)) and not (layer1_outputs(4675));
    layer2_outputs(8852) <= (layer1_outputs(3215)) and (layer1_outputs(264));
    layer2_outputs(8853) <= not(layer1_outputs(7426));
    layer2_outputs(8854) <= not(layer1_outputs(9845));
    layer2_outputs(8855) <= (layer1_outputs(8521)) or (layer1_outputs(8405));
    layer2_outputs(8856) <= layer1_outputs(8049);
    layer2_outputs(8857) <= not(layer1_outputs(9300));
    layer2_outputs(8858) <= (layer1_outputs(992)) and not (layer1_outputs(550));
    layer2_outputs(8859) <= layer1_outputs(8299);
    layer2_outputs(8860) <= not(layer1_outputs(1238));
    layer2_outputs(8861) <= not((layer1_outputs(1866)) xor (layer1_outputs(1699)));
    layer2_outputs(8862) <= not(layer1_outputs(5888)) or (layer1_outputs(8067));
    layer2_outputs(8863) <= not((layer1_outputs(3368)) xor (layer1_outputs(8149)));
    layer2_outputs(8864) <= (layer1_outputs(4512)) or (layer1_outputs(3219));
    layer2_outputs(8865) <= not(layer1_outputs(9561));
    layer2_outputs(8866) <= layer1_outputs(9408);
    layer2_outputs(8867) <= not((layer1_outputs(8071)) and (layer1_outputs(5561)));
    layer2_outputs(8868) <= not(layer1_outputs(2784));
    layer2_outputs(8869) <= layer1_outputs(3407);
    layer2_outputs(8870) <= not(layer1_outputs(4605)) or (layer1_outputs(6660));
    layer2_outputs(8871) <= (layer1_outputs(10200)) and not (layer1_outputs(5017));
    layer2_outputs(8872) <= '0';
    layer2_outputs(8873) <= (layer1_outputs(8305)) and not (layer1_outputs(8976));
    layer2_outputs(8874) <= (layer1_outputs(9092)) xor (layer1_outputs(4921));
    layer2_outputs(8875) <= layer1_outputs(4154);
    layer2_outputs(8876) <= not(layer1_outputs(2188));
    layer2_outputs(8877) <= not((layer1_outputs(4449)) xor (layer1_outputs(8509)));
    layer2_outputs(8878) <= not((layer1_outputs(4697)) xor (layer1_outputs(417)));
    layer2_outputs(8879) <= (layer1_outputs(8948)) and not (layer1_outputs(4393));
    layer2_outputs(8880) <= layer1_outputs(7815);
    layer2_outputs(8881) <= not((layer1_outputs(47)) or (layer1_outputs(8348)));
    layer2_outputs(8882) <= (layer1_outputs(9889)) or (layer1_outputs(2409));
    layer2_outputs(8883) <= not((layer1_outputs(803)) and (layer1_outputs(7475)));
    layer2_outputs(8884) <= (layer1_outputs(4004)) and not (layer1_outputs(4813));
    layer2_outputs(8885) <= not(layer1_outputs(6650));
    layer2_outputs(8886) <= not((layer1_outputs(1118)) or (layer1_outputs(347)));
    layer2_outputs(8887) <= layer1_outputs(7778);
    layer2_outputs(8888) <= layer1_outputs(4532);
    layer2_outputs(8889) <= not(layer1_outputs(9599));
    layer2_outputs(8890) <= not((layer1_outputs(3888)) and (layer1_outputs(9196)));
    layer2_outputs(8891) <= not(layer1_outputs(2150));
    layer2_outputs(8892) <= not(layer1_outputs(1059)) or (layer1_outputs(6693));
    layer2_outputs(8893) <= layer1_outputs(1067);
    layer2_outputs(8894) <= not(layer1_outputs(2080));
    layer2_outputs(8895) <= (layer1_outputs(8663)) xor (layer1_outputs(7100));
    layer2_outputs(8896) <= (layer1_outputs(4263)) xor (layer1_outputs(8896));
    layer2_outputs(8897) <= not(layer1_outputs(4525));
    layer2_outputs(8898) <= not((layer1_outputs(9136)) and (layer1_outputs(9865)));
    layer2_outputs(8899) <= layer1_outputs(3780);
    layer2_outputs(8900) <= not(layer1_outputs(9779)) or (layer1_outputs(7649));
    layer2_outputs(8901) <= (layer1_outputs(3882)) xor (layer1_outputs(6969));
    layer2_outputs(8902) <= (layer1_outputs(8145)) xor (layer1_outputs(10184));
    layer2_outputs(8903) <= not(layer1_outputs(2835));
    layer2_outputs(8904) <= not((layer1_outputs(9556)) xor (layer1_outputs(4766)));
    layer2_outputs(8905) <= not((layer1_outputs(8997)) xor (layer1_outputs(4434)));
    layer2_outputs(8906) <= layer1_outputs(4194);
    layer2_outputs(8907) <= (layer1_outputs(7512)) and not (layer1_outputs(9952));
    layer2_outputs(8908) <= not(layer1_outputs(8680)) or (layer1_outputs(675));
    layer2_outputs(8909) <= not(layer1_outputs(1939));
    layer2_outputs(8910) <= not(layer1_outputs(8286));
    layer2_outputs(8911) <= layer1_outputs(2479);
    layer2_outputs(8912) <= not((layer1_outputs(5297)) and (layer1_outputs(3012)));
    layer2_outputs(8913) <= layer1_outputs(1864);
    layer2_outputs(8914) <= not(layer1_outputs(7760)) or (layer1_outputs(4665));
    layer2_outputs(8915) <= (layer1_outputs(603)) and (layer1_outputs(7220));
    layer2_outputs(8916) <= (layer1_outputs(9425)) or (layer1_outputs(1324));
    layer2_outputs(8917) <= (layer1_outputs(1066)) and not (layer1_outputs(3834));
    layer2_outputs(8918) <= not(layer1_outputs(9427));
    layer2_outputs(8919) <= (layer1_outputs(398)) xor (layer1_outputs(2933));
    layer2_outputs(8920) <= (layer1_outputs(1973)) and not (layer1_outputs(3044));
    layer2_outputs(8921) <= layer1_outputs(8437);
    layer2_outputs(8922) <= layer1_outputs(3802);
    layer2_outputs(8923) <= layer1_outputs(4098);
    layer2_outputs(8924) <= layer1_outputs(9507);
    layer2_outputs(8925) <= (layer1_outputs(1681)) and not (layer1_outputs(1053));
    layer2_outputs(8926) <= not(layer1_outputs(6329));
    layer2_outputs(8927) <= not(layer1_outputs(6193));
    layer2_outputs(8928) <= (layer1_outputs(6315)) or (layer1_outputs(5063));
    layer2_outputs(8929) <= not(layer1_outputs(8166));
    layer2_outputs(8930) <= not((layer1_outputs(333)) xor (layer1_outputs(4881)));
    layer2_outputs(8931) <= layer1_outputs(2309);
    layer2_outputs(8932) <= not((layer1_outputs(6360)) and (layer1_outputs(8860)));
    layer2_outputs(8933) <= not(layer1_outputs(117));
    layer2_outputs(8934) <= not((layer1_outputs(7542)) xor (layer1_outputs(2592)));
    layer2_outputs(8935) <= not((layer1_outputs(8675)) xor (layer1_outputs(6792)));
    layer2_outputs(8936) <= (layer1_outputs(8135)) and not (layer1_outputs(5936));
    layer2_outputs(8937) <= (layer1_outputs(913)) xor (layer1_outputs(4289));
    layer2_outputs(8938) <= not(layer1_outputs(10201)) or (layer1_outputs(3897));
    layer2_outputs(8939) <= not(layer1_outputs(2122));
    layer2_outputs(8940) <= layer1_outputs(5672);
    layer2_outputs(8941) <= not(layer1_outputs(2546)) or (layer1_outputs(10151));
    layer2_outputs(8942) <= not(layer1_outputs(9751)) or (layer1_outputs(1638));
    layer2_outputs(8943) <= not(layer1_outputs(3091));
    layer2_outputs(8944) <= layer1_outputs(5786);
    layer2_outputs(8945) <= not((layer1_outputs(9704)) xor (layer1_outputs(16)));
    layer2_outputs(8946) <= layer1_outputs(7120);
    layer2_outputs(8947) <= not(layer1_outputs(4158));
    layer2_outputs(8948) <= layer1_outputs(7414);
    layer2_outputs(8949) <= not((layer1_outputs(837)) xor (layer1_outputs(786)));
    layer2_outputs(8950) <= not(layer1_outputs(641));
    layer2_outputs(8951) <= layer1_outputs(144);
    layer2_outputs(8952) <= not((layer1_outputs(3722)) xor (layer1_outputs(7131)));
    layer2_outputs(8953) <= layer1_outputs(4739);
    layer2_outputs(8954) <= not(layer1_outputs(8581));
    layer2_outputs(8955) <= (layer1_outputs(1616)) or (layer1_outputs(2351));
    layer2_outputs(8956) <= not(layer1_outputs(5808));
    layer2_outputs(8957) <= not(layer1_outputs(6720)) or (layer1_outputs(315));
    layer2_outputs(8958) <= (layer1_outputs(4699)) xor (layer1_outputs(7991));
    layer2_outputs(8959) <= layer1_outputs(1013);
    layer2_outputs(8960) <= layer1_outputs(440);
    layer2_outputs(8961) <= not(layer1_outputs(5678));
    layer2_outputs(8962) <= layer1_outputs(3392);
    layer2_outputs(8963) <= not(layer1_outputs(6229));
    layer2_outputs(8964) <= not((layer1_outputs(6526)) or (layer1_outputs(379)));
    layer2_outputs(8965) <= (layer1_outputs(8622)) xor (layer1_outputs(9448));
    layer2_outputs(8966) <= not(layer1_outputs(7265));
    layer2_outputs(8967) <= (layer1_outputs(6374)) xor (layer1_outputs(106));
    layer2_outputs(8968) <= not((layer1_outputs(3615)) and (layer1_outputs(4571)));
    layer2_outputs(8969) <= (layer1_outputs(6311)) and (layer1_outputs(4399));
    layer2_outputs(8970) <= (layer1_outputs(1559)) or (layer1_outputs(3414));
    layer2_outputs(8971) <= not(layer1_outputs(8081));
    layer2_outputs(8972) <= not(layer1_outputs(3864)) or (layer1_outputs(4771));
    layer2_outputs(8973) <= not(layer1_outputs(4324));
    layer2_outputs(8974) <= layer1_outputs(2259);
    layer2_outputs(8975) <= not(layer1_outputs(1953));
    layer2_outputs(8976) <= not((layer1_outputs(4062)) xor (layer1_outputs(9440)));
    layer2_outputs(8977) <= not(layer1_outputs(4266));
    layer2_outputs(8978) <= (layer1_outputs(6911)) and not (layer1_outputs(2299));
    layer2_outputs(8979) <= not((layer1_outputs(2547)) and (layer1_outputs(7989)));
    layer2_outputs(8980) <= not((layer1_outputs(3123)) xor (layer1_outputs(4949)));
    layer2_outputs(8981) <= layer1_outputs(8469);
    layer2_outputs(8982) <= layer1_outputs(4220);
    layer2_outputs(8983) <= layer1_outputs(9637);
    layer2_outputs(8984) <= not(layer1_outputs(8254)) or (layer1_outputs(9125));
    layer2_outputs(8985) <= layer1_outputs(3865);
    layer2_outputs(8986) <= (layer1_outputs(574)) and not (layer1_outputs(3659));
    layer2_outputs(8987) <= not(layer1_outputs(2666));
    layer2_outputs(8988) <= not(layer1_outputs(3076)) or (layer1_outputs(6593));
    layer2_outputs(8989) <= not((layer1_outputs(710)) or (layer1_outputs(9369)));
    layer2_outputs(8990) <= not((layer1_outputs(3742)) xor (layer1_outputs(3353)));
    layer2_outputs(8991) <= not((layer1_outputs(1055)) or (layer1_outputs(3511)));
    layer2_outputs(8992) <= layer1_outputs(3006);
    layer2_outputs(8993) <= not(layer1_outputs(5333));
    layer2_outputs(8994) <= not((layer1_outputs(8998)) and (layer1_outputs(5859)));
    layer2_outputs(8995) <= (layer1_outputs(6419)) and not (layer1_outputs(1095));
    layer2_outputs(8996) <= layer1_outputs(5074);
    layer2_outputs(8997) <= not((layer1_outputs(874)) and (layer1_outputs(6450)));
    layer2_outputs(8998) <= not(layer1_outputs(1169));
    layer2_outputs(8999) <= not(layer1_outputs(5182));
    layer2_outputs(9000) <= layer1_outputs(2337);
    layer2_outputs(9001) <= '1';
    layer2_outputs(9002) <= (layer1_outputs(9703)) and not (layer1_outputs(3304));
    layer2_outputs(9003) <= layer1_outputs(5367);
    layer2_outputs(9004) <= not(layer1_outputs(1707));
    layer2_outputs(9005) <= (layer1_outputs(1768)) and (layer1_outputs(885));
    layer2_outputs(9006) <= not((layer1_outputs(1592)) xor (layer1_outputs(5868)));
    layer2_outputs(9007) <= layer1_outputs(8089);
    layer2_outputs(9008) <= not(layer1_outputs(4973)) or (layer1_outputs(5310));
    layer2_outputs(9009) <= '0';
    layer2_outputs(9010) <= not(layer1_outputs(2062));
    layer2_outputs(9011) <= (layer1_outputs(2130)) xor (layer1_outputs(5465));
    layer2_outputs(9012) <= not(layer1_outputs(9560));
    layer2_outputs(9013) <= layer1_outputs(1109);
    layer2_outputs(9014) <= not(layer1_outputs(4179)) or (layer1_outputs(7634));
    layer2_outputs(9015) <= (layer1_outputs(6542)) and not (layer1_outputs(1632));
    layer2_outputs(9016) <= not((layer1_outputs(3456)) xor (layer1_outputs(6406)));
    layer2_outputs(9017) <= not((layer1_outputs(6985)) xor (layer1_outputs(253)));
    layer2_outputs(9018) <= not(layer1_outputs(338));
    layer2_outputs(9019) <= (layer1_outputs(5737)) and (layer1_outputs(7481));
    layer2_outputs(9020) <= (layer1_outputs(3289)) or (layer1_outputs(4556));
    layer2_outputs(9021) <= (layer1_outputs(8009)) xor (layer1_outputs(6120));
    layer2_outputs(9022) <= (layer1_outputs(9653)) xor (layer1_outputs(1756));
    layer2_outputs(9023) <= layer1_outputs(1674);
    layer2_outputs(9024) <= not(layer1_outputs(1819)) or (layer1_outputs(2535));
    layer2_outputs(9025) <= not(layer1_outputs(9433));
    layer2_outputs(9026) <= not(layer1_outputs(3491));
    layer2_outputs(9027) <= (layer1_outputs(7064)) or (layer1_outputs(9790));
    layer2_outputs(9028) <= layer1_outputs(4855);
    layer2_outputs(9029) <= not((layer1_outputs(2510)) and (layer1_outputs(10234)));
    layer2_outputs(9030) <= (layer1_outputs(7809)) and (layer1_outputs(1798));
    layer2_outputs(9031) <= not(layer1_outputs(7220));
    layer2_outputs(9032) <= layer1_outputs(5754);
    layer2_outputs(9033) <= not((layer1_outputs(6103)) xor (layer1_outputs(8787)));
    layer2_outputs(9034) <= not(layer1_outputs(1785));
    layer2_outputs(9035) <= layer1_outputs(191);
    layer2_outputs(9036) <= not(layer1_outputs(8926));
    layer2_outputs(9037) <= not(layer1_outputs(960));
    layer2_outputs(9038) <= (layer1_outputs(6165)) and (layer1_outputs(1888));
    layer2_outputs(9039) <= not((layer1_outputs(7574)) xor (layer1_outputs(504)));
    layer2_outputs(9040) <= not(layer1_outputs(4942));
    layer2_outputs(9041) <= layer1_outputs(7818);
    layer2_outputs(9042) <= (layer1_outputs(5653)) and not (layer1_outputs(5307));
    layer2_outputs(9043) <= (layer1_outputs(6989)) and not (layer1_outputs(3358));
    layer2_outputs(9044) <= not(layer1_outputs(7903));
    layer2_outputs(9045) <= layer1_outputs(2925);
    layer2_outputs(9046) <= (layer1_outputs(4211)) or (layer1_outputs(7885));
    layer2_outputs(9047) <= (layer1_outputs(2738)) xor (layer1_outputs(1052));
    layer2_outputs(9048) <= layer1_outputs(5388);
    layer2_outputs(9049) <= layer1_outputs(3791);
    layer2_outputs(9050) <= layer1_outputs(7142);
    layer2_outputs(9051) <= not(layer1_outputs(10038)) or (layer1_outputs(8338));
    layer2_outputs(9052) <= (layer1_outputs(3609)) and (layer1_outputs(3766));
    layer2_outputs(9053) <= not((layer1_outputs(5283)) or (layer1_outputs(6324)));
    layer2_outputs(9054) <= layer1_outputs(524);
    layer2_outputs(9055) <= not(layer1_outputs(1967));
    layer2_outputs(9056) <= (layer1_outputs(9920)) and not (layer1_outputs(7136));
    layer2_outputs(9057) <= (layer1_outputs(8232)) and not (layer1_outputs(762));
    layer2_outputs(9058) <= layer1_outputs(4575);
    layer2_outputs(9059) <= not(layer1_outputs(459)) or (layer1_outputs(6215));
    layer2_outputs(9060) <= not(layer1_outputs(9622)) or (layer1_outputs(8044));
    layer2_outputs(9061) <= layer1_outputs(7469);
    layer2_outputs(9062) <= (layer1_outputs(4074)) and not (layer1_outputs(9566));
    layer2_outputs(9063) <= (layer1_outputs(9768)) or (layer1_outputs(9978));
    layer2_outputs(9064) <= (layer1_outputs(7165)) xor (layer1_outputs(1075));
    layer2_outputs(9065) <= (layer1_outputs(5013)) xor (layer1_outputs(6355));
    layer2_outputs(9066) <= not(layer1_outputs(7598));
    layer2_outputs(9067) <= not(layer1_outputs(10229)) or (layer1_outputs(5802));
    layer2_outputs(9068) <= not((layer1_outputs(6847)) or (layer1_outputs(4222)));
    layer2_outputs(9069) <= not(layer1_outputs(2215));
    layer2_outputs(9070) <= '1';
    layer2_outputs(9071) <= not(layer1_outputs(4471));
    layer2_outputs(9072) <= layer1_outputs(7793);
    layer2_outputs(9073) <= not(layer1_outputs(6321));
    layer2_outputs(9074) <= layer1_outputs(9800);
    layer2_outputs(9075) <= not((layer1_outputs(5794)) and (layer1_outputs(297)));
    layer2_outputs(9076) <= not(layer1_outputs(3002));
    layer2_outputs(9077) <= layer1_outputs(1190);
    layer2_outputs(9078) <= layer1_outputs(8450);
    layer2_outputs(9079) <= not(layer1_outputs(1165)) or (layer1_outputs(5564));
    layer2_outputs(9080) <= layer1_outputs(1518);
    layer2_outputs(9081) <= (layer1_outputs(9065)) or (layer1_outputs(8284));
    layer2_outputs(9082) <= (layer1_outputs(9006)) and not (layer1_outputs(2321));
    layer2_outputs(9083) <= layer1_outputs(6866);
    layer2_outputs(9084) <= not((layer1_outputs(3674)) xor (layer1_outputs(1340)));
    layer2_outputs(9085) <= (layer1_outputs(7273)) and not (layer1_outputs(4235));
    layer2_outputs(9086) <= not(layer1_outputs(4407));
    layer2_outputs(9087) <= not(layer1_outputs(9892));
    layer2_outputs(9088) <= not((layer1_outputs(5635)) and (layer1_outputs(3960)));
    layer2_outputs(9089) <= layer1_outputs(9565);
    layer2_outputs(9090) <= (layer1_outputs(475)) and not (layer1_outputs(8184));
    layer2_outputs(9091) <= not(layer1_outputs(3797)) or (layer1_outputs(8454));
    layer2_outputs(9092) <= layer1_outputs(246);
    layer2_outputs(9093) <= layer1_outputs(7503);
    layer2_outputs(9094) <= (layer1_outputs(7795)) or (layer1_outputs(7327));
    layer2_outputs(9095) <= layer1_outputs(291);
    layer2_outputs(9096) <= layer1_outputs(3634);
    layer2_outputs(9097) <= layer1_outputs(86);
    layer2_outputs(9098) <= not((layer1_outputs(4378)) and (layer1_outputs(5826)));
    layer2_outputs(9099) <= (layer1_outputs(5309)) xor (layer1_outputs(1114));
    layer2_outputs(9100) <= not(layer1_outputs(612)) or (layer1_outputs(752));
    layer2_outputs(9101) <= not((layer1_outputs(9301)) or (layer1_outputs(4415)));
    layer2_outputs(9102) <= (layer1_outputs(3635)) or (layer1_outputs(4480));
    layer2_outputs(9103) <= (layer1_outputs(7717)) or (layer1_outputs(1411));
    layer2_outputs(9104) <= (layer1_outputs(7607)) and not (layer1_outputs(1509));
    layer2_outputs(9105) <= not((layer1_outputs(635)) xor (layer1_outputs(9499)));
    layer2_outputs(9106) <= not(layer1_outputs(978)) or (layer1_outputs(9881));
    layer2_outputs(9107) <= (layer1_outputs(9372)) and not (layer1_outputs(7705));
    layer2_outputs(9108) <= not(layer1_outputs(74)) or (layer1_outputs(110));
    layer2_outputs(9109) <= (layer1_outputs(4689)) xor (layer1_outputs(5185));
    layer2_outputs(9110) <= not(layer1_outputs(8654)) or (layer1_outputs(2536));
    layer2_outputs(9111) <= not(layer1_outputs(1220));
    layer2_outputs(9112) <= (layer1_outputs(4670)) xor (layer1_outputs(1904));
    layer2_outputs(9113) <= not(layer1_outputs(3022));
    layer2_outputs(9114) <= not((layer1_outputs(2693)) xor (layer1_outputs(4640)));
    layer2_outputs(9115) <= (layer1_outputs(9597)) and not (layer1_outputs(8));
    layer2_outputs(9116) <= (layer1_outputs(4455)) or (layer1_outputs(8289));
    layer2_outputs(9117) <= not((layer1_outputs(1825)) or (layer1_outputs(443)));
    layer2_outputs(9118) <= not(layer1_outputs(4037)) or (layer1_outputs(1750));
    layer2_outputs(9119) <= layer1_outputs(8628);
    layer2_outputs(9120) <= layer1_outputs(5436);
    layer2_outputs(9121) <= not(layer1_outputs(6749));
    layer2_outputs(9122) <= not((layer1_outputs(4053)) and (layer1_outputs(1931)));
    layer2_outputs(9123) <= layer1_outputs(1248);
    layer2_outputs(9124) <= not((layer1_outputs(2000)) and (layer1_outputs(7330)));
    layer2_outputs(9125) <= (layer1_outputs(7976)) or (layer1_outputs(9861));
    layer2_outputs(9126) <= (layer1_outputs(181)) xor (layer1_outputs(4799));
    layer2_outputs(9127) <= not((layer1_outputs(5858)) or (layer1_outputs(5911)));
    layer2_outputs(9128) <= not((layer1_outputs(7259)) xor (layer1_outputs(1608)));
    layer2_outputs(9129) <= not(layer1_outputs(1507));
    layer2_outputs(9130) <= layer1_outputs(328);
    layer2_outputs(9131) <= (layer1_outputs(611)) or (layer1_outputs(8953));
    layer2_outputs(9132) <= layer1_outputs(6987);
    layer2_outputs(9133) <= layer1_outputs(5658);
    layer2_outputs(9134) <= (layer1_outputs(2908)) xor (layer1_outputs(9409));
    layer2_outputs(9135) <= not((layer1_outputs(7649)) or (layer1_outputs(8708)));
    layer2_outputs(9136) <= layer1_outputs(9371);
    layer2_outputs(9137) <= (layer1_outputs(4487)) xor (layer1_outputs(10056));
    layer2_outputs(9138) <= (layer1_outputs(9870)) or (layer1_outputs(6942));
    layer2_outputs(9139) <= not((layer1_outputs(3486)) and (layer1_outputs(632)));
    layer2_outputs(9140) <= layer1_outputs(4632);
    layer2_outputs(9141) <= layer1_outputs(1037);
    layer2_outputs(9142) <= (layer1_outputs(7583)) and not (layer1_outputs(3753));
    layer2_outputs(9143) <= not(layer1_outputs(6603));
    layer2_outputs(9144) <= not(layer1_outputs(8530)) or (layer1_outputs(2262));
    layer2_outputs(9145) <= layer1_outputs(7640);
    layer2_outputs(9146) <= layer1_outputs(1033);
    layer2_outputs(9147) <= not((layer1_outputs(4300)) and (layer1_outputs(2668)));
    layer2_outputs(9148) <= layer1_outputs(1791);
    layer2_outputs(9149) <= (layer1_outputs(8463)) and not (layer1_outputs(6841));
    layer2_outputs(9150) <= layer1_outputs(906);
    layer2_outputs(9151) <= not(layer1_outputs(6768));
    layer2_outputs(9152) <= (layer1_outputs(8995)) or (layer1_outputs(2045));
    layer2_outputs(9153) <= (layer1_outputs(2214)) xor (layer1_outputs(5553));
    layer2_outputs(9154) <= (layer1_outputs(5913)) and not (layer1_outputs(1578));
    layer2_outputs(9155) <= not((layer1_outputs(8400)) and (layer1_outputs(739)));
    layer2_outputs(9156) <= not(layer1_outputs(5173));
    layer2_outputs(9157) <= not(layer1_outputs(410)) or (layer1_outputs(1122));
    layer2_outputs(9158) <= (layer1_outputs(1068)) xor (layer1_outputs(7683));
    layer2_outputs(9159) <= (layer1_outputs(4042)) or (layer1_outputs(9588));
    layer2_outputs(9160) <= layer1_outputs(6050);
    layer2_outputs(9161) <= (layer1_outputs(926)) and not (layer1_outputs(26));
    layer2_outputs(9162) <= layer1_outputs(8068);
    layer2_outputs(9163) <= not((layer1_outputs(10144)) or (layer1_outputs(7774)));
    layer2_outputs(9164) <= (layer1_outputs(9738)) and not (layer1_outputs(7160));
    layer2_outputs(9165) <= layer1_outputs(2295);
    layer2_outputs(9166) <= not(layer1_outputs(6821)) or (layer1_outputs(600));
    layer2_outputs(9167) <= not(layer1_outputs(923));
    layer2_outputs(9168) <= layer1_outputs(3105);
    layer2_outputs(9169) <= (layer1_outputs(5402)) and not (layer1_outputs(3038));
    layer2_outputs(9170) <= (layer1_outputs(2658)) and not (layer1_outputs(3799));
    layer2_outputs(9171) <= layer1_outputs(1209);
    layer2_outputs(9172) <= layer1_outputs(5375);
    layer2_outputs(9173) <= (layer1_outputs(2115)) xor (layer1_outputs(7532));
    layer2_outputs(9174) <= (layer1_outputs(7380)) and not (layer1_outputs(9402));
    layer2_outputs(9175) <= (layer1_outputs(4515)) xor (layer1_outputs(463));
    layer2_outputs(9176) <= not(layer1_outputs(9522));
    layer2_outputs(9177) <= not(layer1_outputs(5498));
    layer2_outputs(9178) <= (layer1_outputs(1268)) and not (layer1_outputs(4812));
    layer2_outputs(9179) <= layer1_outputs(3047);
    layer2_outputs(9180) <= not(layer1_outputs(9907));
    layer2_outputs(9181) <= (layer1_outputs(9997)) and not (layer1_outputs(8124));
    layer2_outputs(9182) <= layer1_outputs(1704);
    layer2_outputs(9183) <= (layer1_outputs(5831)) xor (layer1_outputs(7427));
    layer2_outputs(9184) <= (layer1_outputs(4033)) and not (layer1_outputs(4923));
    layer2_outputs(9185) <= (layer1_outputs(3415)) xor (layer1_outputs(124));
    layer2_outputs(9186) <= not(layer1_outputs(1511));
    layer2_outputs(9187) <= not((layer1_outputs(7690)) or (layer1_outputs(6223)));
    layer2_outputs(9188) <= not(layer1_outputs(5011)) or (layer1_outputs(4610));
    layer2_outputs(9189) <= not((layer1_outputs(2621)) and (layer1_outputs(7907)));
    layer2_outputs(9190) <= layer1_outputs(1338);
    layer2_outputs(9191) <= not((layer1_outputs(8425)) or (layer1_outputs(2)));
    layer2_outputs(9192) <= (layer1_outputs(2519)) and (layer1_outputs(1390));
    layer2_outputs(9193) <= (layer1_outputs(7974)) or (layer1_outputs(3126));
    layer2_outputs(9194) <= not(layer1_outputs(9644));
    layer2_outputs(9195) <= not(layer1_outputs(4390)) or (layer1_outputs(1079));
    layer2_outputs(9196) <= not((layer1_outputs(3156)) and (layer1_outputs(2659)));
    layer2_outputs(9197) <= layer1_outputs(1269);
    layer2_outputs(9198) <= not(layer1_outputs(5875));
    layer2_outputs(9199) <= layer1_outputs(580);
    layer2_outputs(9200) <= layer1_outputs(5398);
    layer2_outputs(9201) <= not(layer1_outputs(10069));
    layer2_outputs(9202) <= layer1_outputs(6612);
    layer2_outputs(9203) <= not(layer1_outputs(10058)) or (layer1_outputs(6084));
    layer2_outputs(9204) <= not((layer1_outputs(9838)) xor (layer1_outputs(6893)));
    layer2_outputs(9205) <= not(layer1_outputs(749));
    layer2_outputs(9206) <= not((layer1_outputs(676)) or (layer1_outputs(7440)));
    layer2_outputs(9207) <= not(layer1_outputs(4786)) or (layer1_outputs(4429));
    layer2_outputs(9208) <= not(layer1_outputs(6102)) or (layer1_outputs(5075));
    layer2_outputs(9209) <= not(layer1_outputs(1897)) or (layer1_outputs(6873));
    layer2_outputs(9210) <= (layer1_outputs(172)) and not (layer1_outputs(7474));
    layer2_outputs(9211) <= not((layer1_outputs(1737)) or (layer1_outputs(3863)));
    layer2_outputs(9212) <= layer1_outputs(727);
    layer2_outputs(9213) <= layer1_outputs(147);
    layer2_outputs(9214) <= not((layer1_outputs(1159)) and (layer1_outputs(5846)));
    layer2_outputs(9215) <= not(layer1_outputs(2603));
    layer2_outputs(9216) <= layer1_outputs(8079);
    layer2_outputs(9217) <= (layer1_outputs(3573)) and (layer1_outputs(1774));
    layer2_outputs(9218) <= not(layer1_outputs(1468));
    layer2_outputs(9219) <= not((layer1_outputs(249)) or (layer1_outputs(6095)));
    layer2_outputs(9220) <= not(layer1_outputs(4057));
    layer2_outputs(9221) <= (layer1_outputs(1443)) and not (layer1_outputs(5878));
    layer2_outputs(9222) <= not((layer1_outputs(9177)) or (layer1_outputs(8686)));
    layer2_outputs(9223) <= not(layer1_outputs(3029)) or (layer1_outputs(3318));
    layer2_outputs(9224) <= (layer1_outputs(8057)) and not (layer1_outputs(8681));
    layer2_outputs(9225) <= not(layer1_outputs(9104));
    layer2_outputs(9226) <= '0';
    layer2_outputs(9227) <= not(layer1_outputs(862));
    layer2_outputs(9228) <= (layer1_outputs(7575)) or (layer1_outputs(8080));
    layer2_outputs(9229) <= (layer1_outputs(5885)) and (layer1_outputs(9621));
    layer2_outputs(9230) <= (layer1_outputs(4746)) xor (layer1_outputs(5935));
    layer2_outputs(9231) <= layer1_outputs(6146);
    layer2_outputs(9232) <= (layer1_outputs(6723)) and not (layer1_outputs(6326));
    layer2_outputs(9233) <= (layer1_outputs(9701)) xor (layer1_outputs(5523));
    layer2_outputs(9234) <= not((layer1_outputs(3269)) or (layer1_outputs(6976)));
    layer2_outputs(9235) <= layer1_outputs(6039);
    layer2_outputs(9236) <= (layer1_outputs(3354)) xor (layer1_outputs(4839));
    layer2_outputs(9237) <= not(layer1_outputs(1061)) or (layer1_outputs(6057));
    layer2_outputs(9238) <= not(layer1_outputs(10007));
    layer2_outputs(9239) <= layer1_outputs(7931);
    layer2_outputs(9240) <= (layer1_outputs(5787)) and not (layer1_outputs(5452));
    layer2_outputs(9241) <= layer1_outputs(1898);
    layer2_outputs(9242) <= (layer1_outputs(109)) and not (layer1_outputs(7667));
    layer2_outputs(9243) <= not((layer1_outputs(5381)) and (layer1_outputs(9062)));
    layer2_outputs(9244) <= not(layer1_outputs(789)) or (layer1_outputs(1090));
    layer2_outputs(9245) <= (layer1_outputs(6431)) xor (layer1_outputs(9614));
    layer2_outputs(9246) <= not(layer1_outputs(2294)) or (layer1_outputs(2804));
    layer2_outputs(9247) <= not((layer1_outputs(6532)) xor (layer1_outputs(1915)));
    layer2_outputs(9248) <= not(layer1_outputs(2941));
    layer2_outputs(9249) <= not(layer1_outputs(4691));
    layer2_outputs(9250) <= (layer1_outputs(2428)) xor (layer1_outputs(683));
    layer2_outputs(9251) <= not(layer1_outputs(7343)) or (layer1_outputs(8952));
    layer2_outputs(9252) <= '1';
    layer2_outputs(9253) <= (layer1_outputs(548)) and not (layer1_outputs(3325));
    layer2_outputs(9254) <= not(layer1_outputs(565));
    layer2_outputs(9255) <= (layer1_outputs(6423)) and (layer1_outputs(8819));
    layer2_outputs(9256) <= not(layer1_outputs(2699));
    layer2_outputs(9257) <= not((layer1_outputs(7519)) and (layer1_outputs(4648)));
    layer2_outputs(9258) <= layer1_outputs(5341);
    layer2_outputs(9259) <= layer1_outputs(9853);
    layer2_outputs(9260) <= (layer1_outputs(5261)) and not (layer1_outputs(63));
    layer2_outputs(9261) <= not(layer1_outputs(4248)) or (layer1_outputs(10120));
    layer2_outputs(9262) <= not(layer1_outputs(201)) or (layer1_outputs(909));
    layer2_outputs(9263) <= layer1_outputs(459);
    layer2_outputs(9264) <= (layer1_outputs(4995)) or (layer1_outputs(7533));
    layer2_outputs(9265) <= (layer1_outputs(3709)) xor (layer1_outputs(10123));
    layer2_outputs(9266) <= (layer1_outputs(640)) and not (layer1_outputs(2203));
    layer2_outputs(9267) <= (layer1_outputs(5748)) and not (layer1_outputs(8076));
    layer2_outputs(9268) <= (layer1_outputs(7124)) and not (layer1_outputs(5476));
    layer2_outputs(9269) <= (layer1_outputs(6736)) and (layer1_outputs(7044));
    layer2_outputs(9270) <= not(layer1_outputs(5001)) or (layer1_outputs(363));
    layer2_outputs(9271) <= layer1_outputs(2585);
    layer2_outputs(9272) <= (layer1_outputs(1101)) xor (layer1_outputs(9156));
    layer2_outputs(9273) <= (layer1_outputs(1185)) and not (layer1_outputs(5324));
    layer2_outputs(9274) <= not((layer1_outputs(1354)) or (layer1_outputs(6944)));
    layer2_outputs(9275) <= not(layer1_outputs(1716));
    layer2_outputs(9276) <= layer1_outputs(8729);
    layer2_outputs(9277) <= not(layer1_outputs(2411)) or (layer1_outputs(2985));
    layer2_outputs(9278) <= not(layer1_outputs(1454)) or (layer1_outputs(8898));
    layer2_outputs(9279) <= not(layer1_outputs(578));
    layer2_outputs(9280) <= (layer1_outputs(8851)) xor (layer1_outputs(1527));
    layer2_outputs(9281) <= layer1_outputs(4232);
    layer2_outputs(9282) <= (layer1_outputs(3838)) and not (layer1_outputs(6952));
    layer2_outputs(9283) <= layer1_outputs(4582);
    layer2_outputs(9284) <= not((layer1_outputs(4516)) and (layer1_outputs(7683)));
    layer2_outputs(9285) <= not(layer1_outputs(1747));
    layer2_outputs(9286) <= layer1_outputs(9593);
    layer2_outputs(9287) <= (layer1_outputs(3403)) xor (layer1_outputs(7158));
    layer2_outputs(9288) <= (layer1_outputs(2726)) xor (layer1_outputs(436));
    layer2_outputs(9289) <= not((layer1_outputs(4423)) and (layer1_outputs(2294)));
    layer2_outputs(9290) <= layer1_outputs(5965);
    layer2_outputs(9291) <= layer1_outputs(7615);
    layer2_outputs(9292) <= not((layer1_outputs(7864)) or (layer1_outputs(1230)));
    layer2_outputs(9293) <= not(layer1_outputs(6727)) or (layer1_outputs(7920));
    layer2_outputs(9294) <= layer1_outputs(1109);
    layer2_outputs(9295) <= not(layer1_outputs(7113)) or (layer1_outputs(290));
    layer2_outputs(9296) <= not((layer1_outputs(4500)) or (layer1_outputs(45)));
    layer2_outputs(9297) <= not((layer1_outputs(9659)) and (layer1_outputs(5492)));
    layer2_outputs(9298) <= layer1_outputs(1833);
    layer2_outputs(9299) <= not(layer1_outputs(434));
    layer2_outputs(9300) <= layer1_outputs(9700);
    layer2_outputs(9301) <= not(layer1_outputs(4759));
    layer2_outputs(9302) <= layer1_outputs(3739);
    layer2_outputs(9303) <= not(layer1_outputs(4733));
    layer2_outputs(9304) <= not((layer1_outputs(4479)) or (layer1_outputs(2641)));
    layer2_outputs(9305) <= not(layer1_outputs(8229));
    layer2_outputs(9306) <= (layer1_outputs(2361)) and not (layer1_outputs(8704));
    layer2_outputs(9307) <= not((layer1_outputs(9726)) xor (layer1_outputs(10178)));
    layer2_outputs(9308) <= layer1_outputs(8277);
    layer2_outputs(9309) <= not((layer1_outputs(8784)) and (layer1_outputs(5604)));
    layer2_outputs(9310) <= layer1_outputs(8248);
    layer2_outputs(9311) <= (layer1_outputs(3271)) and not (layer1_outputs(6500));
    layer2_outputs(9312) <= (layer1_outputs(9286)) and (layer1_outputs(1491));
    layer2_outputs(9313) <= not((layer1_outputs(9437)) or (layer1_outputs(3762)));
    layer2_outputs(9314) <= not(layer1_outputs(8685));
    layer2_outputs(9315) <= (layer1_outputs(1259)) xor (layer1_outputs(6588));
    layer2_outputs(9316) <= not(layer1_outputs(1206));
    layer2_outputs(9317) <= not((layer1_outputs(5662)) xor (layer1_outputs(2147)));
    layer2_outputs(9318) <= layer1_outputs(3165);
    layer2_outputs(9319) <= layer1_outputs(531);
    layer2_outputs(9320) <= layer1_outputs(1862);
    layer2_outputs(9321) <= layer1_outputs(6343);
    layer2_outputs(9322) <= layer1_outputs(3732);
    layer2_outputs(9323) <= (layer1_outputs(3485)) or (layer1_outputs(5848));
    layer2_outputs(9324) <= (layer1_outputs(9846)) xor (layer1_outputs(7019));
    layer2_outputs(9325) <= not(layer1_outputs(3166));
    layer2_outputs(9326) <= not(layer1_outputs(2752)) or (layer1_outputs(3877));
    layer2_outputs(9327) <= layer1_outputs(3850);
    layer2_outputs(9328) <= not(layer1_outputs(3515));
    layer2_outputs(9329) <= not(layer1_outputs(6618));
    layer2_outputs(9330) <= layer1_outputs(10066);
    layer2_outputs(9331) <= layer1_outputs(4444);
    layer2_outputs(9332) <= (layer1_outputs(8529)) xor (layer1_outputs(9534));
    layer2_outputs(9333) <= layer1_outputs(3811);
    layer2_outputs(9334) <= layer1_outputs(722);
    layer2_outputs(9335) <= not(layer1_outputs(269));
    layer2_outputs(9336) <= not(layer1_outputs(9664));
    layer2_outputs(9337) <= not(layer1_outputs(3578));
    layer2_outputs(9338) <= (layer1_outputs(10118)) and (layer1_outputs(3161));
    layer2_outputs(9339) <= (layer1_outputs(3117)) and not (layer1_outputs(8403));
    layer2_outputs(9340) <= not(layer1_outputs(9896));
    layer2_outputs(9341) <= layer1_outputs(6159);
    layer2_outputs(9342) <= not((layer1_outputs(7739)) xor (layer1_outputs(1599)));
    layer2_outputs(9343) <= not(layer1_outputs(2805));
    layer2_outputs(9344) <= (layer1_outputs(5845)) or (layer1_outputs(850));
    layer2_outputs(9345) <= not((layer1_outputs(7988)) and (layer1_outputs(6448)));
    layer2_outputs(9346) <= (layer1_outputs(7043)) xor (layer1_outputs(5682));
    layer2_outputs(9347) <= layer1_outputs(6683);
    layer2_outputs(9348) <= not((layer1_outputs(8500)) xor (layer1_outputs(3599)));
    layer2_outputs(9349) <= not((layer1_outputs(7695)) xor (layer1_outputs(8749)));
    layer2_outputs(9350) <= not((layer1_outputs(4809)) and (layer1_outputs(5244)));
    layer2_outputs(9351) <= (layer1_outputs(194)) and not (layer1_outputs(6));
    layer2_outputs(9352) <= not((layer1_outputs(1696)) or (layer1_outputs(8572)));
    layer2_outputs(9353) <= layer1_outputs(9420);
    layer2_outputs(9354) <= not(layer1_outputs(4606));
    layer2_outputs(9355) <= (layer1_outputs(9624)) and not (layer1_outputs(6708));
    layer2_outputs(9356) <= (layer1_outputs(9761)) or (layer1_outputs(4047));
    layer2_outputs(9357) <= layer1_outputs(450);
    layer2_outputs(9358) <= not((layer1_outputs(10029)) xor (layer1_outputs(3172)));
    layer2_outputs(9359) <= (layer1_outputs(9)) and not (layer1_outputs(8133));
    layer2_outputs(9360) <= layer1_outputs(2841);
    layer2_outputs(9361) <= not(layer1_outputs(4423));
    layer2_outputs(9362) <= layer1_outputs(492);
    layer2_outputs(9363) <= not(layer1_outputs(2493));
    layer2_outputs(9364) <= not((layer1_outputs(8354)) xor (layer1_outputs(8523)));
    layer2_outputs(9365) <= layer1_outputs(4616);
    layer2_outputs(9366) <= (layer1_outputs(1513)) xor (layer1_outputs(1302));
    layer2_outputs(9367) <= (layer1_outputs(4589)) and not (layer1_outputs(9381));
    layer2_outputs(9368) <= not((layer1_outputs(1876)) and (layer1_outputs(5528)));
    layer2_outputs(9369) <= not(layer1_outputs(8620)) or (layer1_outputs(2061));
    layer2_outputs(9370) <= not(layer1_outputs(9035));
    layer2_outputs(9371) <= layer1_outputs(2270);
    layer2_outputs(9372) <= (layer1_outputs(1482)) and (layer1_outputs(923));
    layer2_outputs(9373) <= (layer1_outputs(9589)) and (layer1_outputs(6147));
    layer2_outputs(9374) <= layer1_outputs(4584);
    layer2_outputs(9375) <= not(layer1_outputs(7965));
    layer2_outputs(9376) <= layer1_outputs(10198);
    layer2_outputs(9377) <= (layer1_outputs(5214)) xor (layer1_outputs(7328));
    layer2_outputs(9378) <= (layer1_outputs(2509)) and (layer1_outputs(5926));
    layer2_outputs(9379) <= layer1_outputs(8364);
    layer2_outputs(9380) <= layer1_outputs(6754);
    layer2_outputs(9381) <= not((layer1_outputs(4290)) xor (layer1_outputs(6003)));
    layer2_outputs(9382) <= layer1_outputs(8652);
    layer2_outputs(9383) <= not(layer1_outputs(4019)) or (layer1_outputs(5476));
    layer2_outputs(9384) <= not(layer1_outputs(2254));
    layer2_outputs(9385) <= layer1_outputs(4945);
    layer2_outputs(9386) <= not(layer1_outputs(3745));
    layer2_outputs(9387) <= (layer1_outputs(6204)) and not (layer1_outputs(4307));
    layer2_outputs(9388) <= layer1_outputs(10204);
    layer2_outputs(9389) <= not((layer1_outputs(7685)) or (layer1_outputs(1085)));
    layer2_outputs(9390) <= not(layer1_outputs(2313));
    layer2_outputs(9391) <= layer1_outputs(4377);
    layer2_outputs(9392) <= not(layer1_outputs(6643)) or (layer1_outputs(231));
    layer2_outputs(9393) <= layer1_outputs(3070);
    layer2_outputs(9394) <= layer1_outputs(3826);
    layer2_outputs(9395) <= (layer1_outputs(2483)) and (layer1_outputs(7095));
    layer2_outputs(9396) <= not(layer1_outputs(4277)) or (layer1_outputs(9288));
    layer2_outputs(9397) <= not((layer1_outputs(6728)) xor (layer1_outputs(5378)));
    layer2_outputs(9398) <= layer1_outputs(7098);
    layer2_outputs(9399) <= (layer1_outputs(7279)) and not (layer1_outputs(6574));
    layer2_outputs(9400) <= (layer1_outputs(7745)) and not (layer1_outputs(7130));
    layer2_outputs(9401) <= layer1_outputs(5322);
    layer2_outputs(9402) <= (layer1_outputs(3514)) or (layer1_outputs(7384));
    layer2_outputs(9403) <= not(layer1_outputs(8743)) or (layer1_outputs(7149));
    layer2_outputs(9404) <= not(layer1_outputs(5539));
    layer2_outputs(9405) <= (layer1_outputs(3519)) and not (layer1_outputs(5272));
    layer2_outputs(9406) <= not((layer1_outputs(1772)) xor (layer1_outputs(2939)));
    layer2_outputs(9407) <= not(layer1_outputs(7690));
    layer2_outputs(9408) <= not(layer1_outputs(3071)) or (layer1_outputs(5654));
    layer2_outputs(9409) <= (layer1_outputs(5879)) and (layer1_outputs(7441));
    layer2_outputs(9410) <= layer1_outputs(1687);
    layer2_outputs(9411) <= (layer1_outputs(9652)) or (layer1_outputs(2336));
    layer2_outputs(9412) <= not(layer1_outputs(5627)) or (layer1_outputs(1789));
    layer2_outputs(9413) <= not((layer1_outputs(6184)) and (layer1_outputs(7494)));
    layer2_outputs(9414) <= (layer1_outputs(6694)) and not (layer1_outputs(8794));
    layer2_outputs(9415) <= not((layer1_outputs(10039)) and (layer1_outputs(9801)));
    layer2_outputs(9416) <= not((layer1_outputs(8807)) or (layer1_outputs(6717)));
    layer2_outputs(9417) <= not(layer1_outputs(9612));
    layer2_outputs(9418) <= not(layer1_outputs(3773));
    layer2_outputs(9419) <= (layer1_outputs(477)) or (layer1_outputs(10186));
    layer2_outputs(9420) <= (layer1_outputs(7154)) or (layer1_outputs(10036));
    layer2_outputs(9421) <= not(layer1_outputs(982));
    layer2_outputs(9422) <= not((layer1_outputs(252)) and (layer1_outputs(745)));
    layer2_outputs(9423) <= not(layer1_outputs(2883));
    layer2_outputs(9424) <= (layer1_outputs(3212)) xor (layer1_outputs(6075));
    layer2_outputs(9425) <= layer1_outputs(6383);
    layer2_outputs(9426) <= not((layer1_outputs(8328)) or (layer1_outputs(5486)));
    layer2_outputs(9427) <= not(layer1_outputs(5799)) or (layer1_outputs(3790));
    layer2_outputs(9428) <= not(layer1_outputs(8877));
    layer2_outputs(9429) <= not(layer1_outputs(5701));
    layer2_outputs(9430) <= not(layer1_outputs(7983)) or (layer1_outputs(1317));
    layer2_outputs(9431) <= (layer1_outputs(4891)) or (layer1_outputs(7715));
    layer2_outputs(9432) <= not((layer1_outputs(8734)) and (layer1_outputs(7095)));
    layer2_outputs(9433) <= not((layer1_outputs(4892)) or (layer1_outputs(317)));
    layer2_outputs(9434) <= (layer1_outputs(6980)) or (layer1_outputs(2495));
    layer2_outputs(9435) <= not((layer1_outputs(10030)) xor (layer1_outputs(1956)));
    layer2_outputs(9436) <= layer1_outputs(7869);
    layer2_outputs(9437) <= not(layer1_outputs(6966)) or (layer1_outputs(7969));
    layer2_outputs(9438) <= layer1_outputs(2985);
    layer2_outputs(9439) <= not(layer1_outputs(5032)) or (layer1_outputs(6892));
    layer2_outputs(9440) <= (layer1_outputs(8)) or (layer1_outputs(4010));
    layer2_outputs(9441) <= layer1_outputs(8910);
    layer2_outputs(9442) <= (layer1_outputs(3934)) and not (layer1_outputs(9171));
    layer2_outputs(9443) <= not((layer1_outputs(4559)) xor (layer1_outputs(1656)));
    layer2_outputs(9444) <= not(layer1_outputs(1083));
    layer2_outputs(9445) <= not((layer1_outputs(1730)) and (layer1_outputs(9631)));
    layer2_outputs(9446) <= layer1_outputs(171);
    layer2_outputs(9447) <= not((layer1_outputs(5777)) or (layer1_outputs(7425)));
    layer2_outputs(9448) <= layer1_outputs(3662);
    layer2_outputs(9449) <= layer1_outputs(4940);
    layer2_outputs(9450) <= layer1_outputs(1170);
    layer2_outputs(9451) <= layer1_outputs(4966);
    layer2_outputs(9452) <= (layer1_outputs(1044)) and not (layer1_outputs(4103));
    layer2_outputs(9453) <= not(layer1_outputs(9957));
    layer2_outputs(9454) <= not(layer1_outputs(8689)) or (layer1_outputs(7074));
    layer2_outputs(9455) <= layer1_outputs(4208);
    layer2_outputs(9456) <= (layer1_outputs(844)) and (layer1_outputs(1184));
    layer2_outputs(9457) <= not((layer1_outputs(8366)) and (layer1_outputs(9978)));
    layer2_outputs(9458) <= layer1_outputs(5622);
    layer2_outputs(9459) <= layer1_outputs(2442);
    layer2_outputs(9460) <= not(layer1_outputs(1136));
    layer2_outputs(9461) <= (layer1_outputs(96)) xor (layer1_outputs(4654));
    layer2_outputs(9462) <= not(layer1_outputs(374)) or (layer1_outputs(4009));
    layer2_outputs(9463) <= not(layer1_outputs(6413));
    layer2_outputs(9464) <= layer1_outputs(3672);
    layer2_outputs(9465) <= not(layer1_outputs(804));
    layer2_outputs(9466) <= layer1_outputs(3657);
    layer2_outputs(9467) <= not(layer1_outputs(4970));
    layer2_outputs(9468) <= (layer1_outputs(9039)) and not (layer1_outputs(861));
    layer2_outputs(9469) <= '0';
    layer2_outputs(9470) <= layer1_outputs(7769);
    layer2_outputs(9471) <= not((layer1_outputs(1073)) and (layer1_outputs(3360)));
    layer2_outputs(9472) <= layer1_outputs(969);
    layer2_outputs(9473) <= not(layer1_outputs(7972)) or (layer1_outputs(3566));
    layer2_outputs(9474) <= not(layer1_outputs(3486)) or (layer1_outputs(125));
    layer2_outputs(9475) <= not((layer1_outputs(5299)) xor (layer1_outputs(132)));
    layer2_outputs(9476) <= not(layer1_outputs(5211));
    layer2_outputs(9477) <= (layer1_outputs(9134)) xor (layer1_outputs(5807));
    layer2_outputs(9478) <= not(layer1_outputs(4722));
    layer2_outputs(9479) <= layer1_outputs(4401);
    layer2_outputs(9480) <= layer1_outputs(7253);
    layer2_outputs(9481) <= not(layer1_outputs(8319)) or (layer1_outputs(4898));
    layer2_outputs(9482) <= not(layer1_outputs(4941));
    layer2_outputs(9483) <= layer1_outputs(553);
    layer2_outputs(9484) <= not(layer1_outputs(6896));
    layer2_outputs(9485) <= layer1_outputs(8178);
    layer2_outputs(9486) <= not((layer1_outputs(604)) xor (layer1_outputs(8087)));
    layer2_outputs(9487) <= not((layer1_outputs(9444)) xor (layer1_outputs(7092)));
    layer2_outputs(9488) <= not(layer1_outputs(1550)) or (layer1_outputs(7296));
    layer2_outputs(9489) <= not(layer1_outputs(2157));
    layer2_outputs(9490) <= not(layer1_outputs(9466)) or (layer1_outputs(7492));
    layer2_outputs(9491) <= not(layer1_outputs(2035)) or (layer1_outputs(4684));
    layer2_outputs(9492) <= layer1_outputs(6845);
    layer2_outputs(9493) <= not((layer1_outputs(6787)) or (layer1_outputs(3210)));
    layer2_outputs(9494) <= (layer1_outputs(6793)) xor (layer1_outputs(1516));
    layer2_outputs(9495) <= layer1_outputs(10201);
    layer2_outputs(9496) <= (layer1_outputs(4315)) and not (layer1_outputs(2205));
    layer2_outputs(9497) <= not(layer1_outputs(528));
    layer2_outputs(9498) <= not(layer1_outputs(4290)) or (layer1_outputs(3635));
    layer2_outputs(9499) <= layer1_outputs(5280);
    layer2_outputs(9500) <= layer1_outputs(6875);
    layer2_outputs(9501) <= not(layer1_outputs(6589)) or (layer1_outputs(2228));
    layer2_outputs(9502) <= not(layer1_outputs(3793));
    layer2_outputs(9503) <= not((layer1_outputs(9072)) or (layer1_outputs(2526)));
    layer2_outputs(9504) <= not(layer1_outputs(8300));
    layer2_outputs(9505) <= layer1_outputs(4217);
    layer2_outputs(9506) <= not(layer1_outputs(9774));
    layer2_outputs(9507) <= not(layer1_outputs(2273));
    layer2_outputs(9508) <= not((layer1_outputs(2518)) and (layer1_outputs(2388)));
    layer2_outputs(9509) <= not(layer1_outputs(10098)) or (layer1_outputs(8803));
    layer2_outputs(9510) <= (layer1_outputs(9596)) and (layer1_outputs(3084));
    layer2_outputs(9511) <= not((layer1_outputs(8452)) and (layer1_outputs(7128)));
    layer2_outputs(9512) <= (layer1_outputs(1424)) or (layer1_outputs(6777));
    layer2_outputs(9513) <= (layer1_outputs(9112)) and (layer1_outputs(2773));
    layer2_outputs(9514) <= not((layer1_outputs(9269)) xor (layer1_outputs(911)));
    layer2_outputs(9515) <= not(layer1_outputs(2077)) or (layer1_outputs(401));
    layer2_outputs(9516) <= not(layer1_outputs(401));
    layer2_outputs(9517) <= (layer1_outputs(1891)) and not (layer1_outputs(224));
    layer2_outputs(9518) <= not((layer1_outputs(6442)) and (layer1_outputs(3126)));
    layer2_outputs(9519) <= not(layer1_outputs(1734));
    layer2_outputs(9520) <= not(layer1_outputs(6834));
    layer2_outputs(9521) <= layer1_outputs(261);
    layer2_outputs(9522) <= (layer1_outputs(9589)) xor (layer1_outputs(7749));
    layer2_outputs(9523) <= layer1_outputs(4518);
    layer2_outputs(9524) <= layer1_outputs(8768);
    layer2_outputs(9525) <= (layer1_outputs(6611)) and not (layer1_outputs(8396));
    layer2_outputs(9526) <= not((layer1_outputs(6794)) and (layer1_outputs(601)));
    layer2_outputs(9527) <= layer1_outputs(2694);
    layer2_outputs(9528) <= (layer1_outputs(8731)) and not (layer1_outputs(3584));
    layer2_outputs(9529) <= (layer1_outputs(3316)) xor (layer1_outputs(710));
    layer2_outputs(9530) <= layer1_outputs(3215);
    layer2_outputs(9531) <= not(layer1_outputs(9333));
    layer2_outputs(9532) <= layer1_outputs(9832);
    layer2_outputs(9533) <= not((layer1_outputs(6531)) xor (layer1_outputs(2412)));
    layer2_outputs(9534) <= layer1_outputs(537);
    layer2_outputs(9535) <= not(layer1_outputs(7236)) or (layer1_outputs(3888));
    layer2_outputs(9536) <= (layer1_outputs(9234)) and not (layer1_outputs(1782));
    layer2_outputs(9537) <= not((layer1_outputs(7779)) or (layer1_outputs(1198)));
    layer2_outputs(9538) <= not(layer1_outputs(6456));
    layer2_outputs(9539) <= not(layer1_outputs(8841));
    layer2_outputs(9540) <= (layer1_outputs(3665)) and not (layer1_outputs(3353));
    layer2_outputs(9541) <= layer1_outputs(6905);
    layer2_outputs(9542) <= not((layer1_outputs(1017)) or (layer1_outputs(2415)));
    layer2_outputs(9543) <= not(layer1_outputs(6047));
    layer2_outputs(9544) <= not(layer1_outputs(5601));
    layer2_outputs(9545) <= layer1_outputs(6188);
    layer2_outputs(9546) <= layer1_outputs(2814);
    layer2_outputs(9547) <= not((layer1_outputs(1424)) xor (layer1_outputs(6268)));
    layer2_outputs(9548) <= not(layer1_outputs(4991)) or (layer1_outputs(628));
    layer2_outputs(9549) <= layer1_outputs(1422);
    layer2_outputs(9550) <= not(layer1_outputs(4654));
    layer2_outputs(9551) <= not((layer1_outputs(6261)) or (layer1_outputs(6484)));
    layer2_outputs(9552) <= (layer1_outputs(3046)) and not (layer1_outputs(7689));
    layer2_outputs(9553) <= (layer1_outputs(4239)) and not (layer1_outputs(9991));
    layer2_outputs(9554) <= not(layer1_outputs(3674));
    layer2_outputs(9555) <= (layer1_outputs(9358)) xor (layer1_outputs(8360));
    layer2_outputs(9556) <= not(layer1_outputs(3946));
    layer2_outputs(9557) <= not(layer1_outputs(10084));
    layer2_outputs(9558) <= not(layer1_outputs(5352));
    layer2_outputs(9559) <= not(layer1_outputs(2502)) or (layer1_outputs(10146));
    layer2_outputs(9560) <= not(layer1_outputs(4800));
    layer2_outputs(9561) <= layer1_outputs(1693);
    layer2_outputs(9562) <= layer1_outputs(2338);
    layer2_outputs(9563) <= layer1_outputs(8467);
    layer2_outputs(9564) <= (layer1_outputs(4105)) and (layer1_outputs(634));
    layer2_outputs(9565) <= (layer1_outputs(7149)) xor (layer1_outputs(6543));
    layer2_outputs(9566) <= not(layer1_outputs(8081));
    layer2_outputs(9567) <= not((layer1_outputs(6280)) and (layer1_outputs(5900)));
    layer2_outputs(9568) <= not(layer1_outputs(2301));
    layer2_outputs(9569) <= not(layer1_outputs(9707)) or (layer1_outputs(8132));
    layer2_outputs(9570) <= '0';
    layer2_outputs(9571) <= layer1_outputs(7159);
    layer2_outputs(9572) <= not(layer1_outputs(6984)) or (layer1_outputs(8693));
    layer2_outputs(9573) <= (layer1_outputs(1133)) and not (layer1_outputs(2107));
    layer2_outputs(9574) <= layer1_outputs(2797);
    layer2_outputs(9575) <= (layer1_outputs(2383)) xor (layer1_outputs(7307));
    layer2_outputs(9576) <= layer1_outputs(4805);
    layer2_outputs(9577) <= layer1_outputs(2917);
    layer2_outputs(9578) <= layer1_outputs(4963);
    layer2_outputs(9579) <= not(layer1_outputs(7290));
    layer2_outputs(9580) <= not((layer1_outputs(2928)) or (layer1_outputs(3910)));
    layer2_outputs(9581) <= not(layer1_outputs(7377));
    layer2_outputs(9582) <= (layer1_outputs(2581)) xor (layer1_outputs(4406));
    layer2_outputs(9583) <= not((layer1_outputs(4854)) xor (layer1_outputs(8514)));
    layer2_outputs(9584) <= (layer1_outputs(4382)) or (layer1_outputs(7288));
    layer2_outputs(9585) <= (layer1_outputs(2983)) and not (layer1_outputs(1300));
    layer2_outputs(9586) <= (layer1_outputs(9450)) xor (layer1_outputs(4002));
    layer2_outputs(9587) <= not((layer1_outputs(821)) and (layer1_outputs(3389)));
    layer2_outputs(9588) <= not(layer1_outputs(6260)) or (layer1_outputs(5530));
    layer2_outputs(9589) <= (layer1_outputs(71)) or (layer1_outputs(5710));
    layer2_outputs(9590) <= layer1_outputs(3918);
    layer2_outputs(9591) <= not(layer1_outputs(2648)) or (layer1_outputs(7979));
    layer2_outputs(9592) <= layer1_outputs(3555);
    layer2_outputs(9593) <= not(layer1_outputs(8964));
    layer2_outputs(9594) <= not(layer1_outputs(2793));
    layer2_outputs(9595) <= not((layer1_outputs(8138)) or (layer1_outputs(6713)));
    layer2_outputs(9596) <= layer1_outputs(5127);
    layer2_outputs(9597) <= not(layer1_outputs(8578)) or (layer1_outputs(2413));
    layer2_outputs(9598) <= (layer1_outputs(2836)) and not (layer1_outputs(4133));
    layer2_outputs(9599) <= layer1_outputs(2278);
    layer2_outputs(9600) <= layer1_outputs(5538);
    layer2_outputs(9601) <= (layer1_outputs(670)) and not (layer1_outputs(1575));
    layer2_outputs(9602) <= not((layer1_outputs(3565)) xor (layer1_outputs(6203)));
    layer2_outputs(9603) <= (layer1_outputs(5410)) xor (layer1_outputs(2897));
    layer2_outputs(9604) <= (layer1_outputs(8162)) and not (layer1_outputs(5383));
    layer2_outputs(9605) <= (layer1_outputs(8353)) and not (layer1_outputs(4714));
    layer2_outputs(9606) <= not(layer1_outputs(966));
    layer2_outputs(9607) <= (layer1_outputs(8894)) and not (layer1_outputs(7126));
    layer2_outputs(9608) <= '0';
    layer2_outputs(9609) <= not(layer1_outputs(8310));
    layer2_outputs(9610) <= (layer1_outputs(1031)) xor (layer1_outputs(7953));
    layer2_outputs(9611) <= not(layer1_outputs(6027));
    layer2_outputs(9612) <= layer1_outputs(4847);
    layer2_outputs(9613) <= layer1_outputs(8218);
    layer2_outputs(9614) <= not((layer1_outputs(2154)) or (layer1_outputs(5050)));
    layer2_outputs(9615) <= not(layer1_outputs(5845));
    layer2_outputs(9616) <= not((layer1_outputs(7074)) xor (layer1_outputs(5941)));
    layer2_outputs(9617) <= layer1_outputs(9606);
    layer2_outputs(9618) <= not(layer1_outputs(6981));
    layer2_outputs(9619) <= (layer1_outputs(2465)) xor (layer1_outputs(2593));
    layer2_outputs(9620) <= layer1_outputs(5864);
    layer2_outputs(9621) <= layer1_outputs(2472);
    layer2_outputs(9622) <= not((layer1_outputs(6516)) and (layer1_outputs(2028)));
    layer2_outputs(9623) <= layer1_outputs(5576);
    layer2_outputs(9624) <= not(layer1_outputs(6110));
    layer2_outputs(9625) <= not(layer1_outputs(8249));
    layer2_outputs(9626) <= '1';
    layer2_outputs(9627) <= not(layer1_outputs(4748)) or (layer1_outputs(747));
    layer2_outputs(9628) <= layer1_outputs(2356);
    layer2_outputs(9629) <= not((layer1_outputs(8064)) or (layer1_outputs(2677)));
    layer2_outputs(9630) <= not((layer1_outputs(5003)) xor (layer1_outputs(4009)));
    layer2_outputs(9631) <= not((layer1_outputs(2182)) and (layer1_outputs(6553)));
    layer2_outputs(9632) <= not((layer1_outputs(1701)) or (layer1_outputs(9082)));
    layer2_outputs(9633) <= not(layer1_outputs(1962));
    layer2_outputs(9634) <= not(layer1_outputs(1828));
    layer2_outputs(9635) <= layer1_outputs(1993);
    layer2_outputs(9636) <= not(layer1_outputs(8891));
    layer2_outputs(9637) <= not(layer1_outputs(6660));
    layer2_outputs(9638) <= (layer1_outputs(5838)) xor (layer1_outputs(3667));
    layer2_outputs(9639) <= not(layer1_outputs(4336)) or (layer1_outputs(9378));
    layer2_outputs(9640) <= not((layer1_outputs(9976)) or (layer1_outputs(8983)));
    layer2_outputs(9641) <= (layer1_outputs(1419)) and (layer1_outputs(8408));
    layer2_outputs(9642) <= not(layer1_outputs(2255));
    layer2_outputs(9643) <= not((layer1_outputs(2999)) or (layer1_outputs(10051)));
    layer2_outputs(9644) <= layer1_outputs(284);
    layer2_outputs(9645) <= (layer1_outputs(6521)) xor (layer1_outputs(5749));
    layer2_outputs(9646) <= not(layer1_outputs(3211));
    layer2_outputs(9647) <= (layer1_outputs(7302)) xor (layer1_outputs(5129));
    layer2_outputs(9648) <= not(layer1_outputs(5027));
    layer2_outputs(9649) <= (layer1_outputs(1184)) or (layer1_outputs(5343));
    layer2_outputs(9650) <= not(layer1_outputs(4604)) or (layer1_outputs(4489));
    layer2_outputs(9651) <= layer1_outputs(6790);
    layer2_outputs(9652) <= layer1_outputs(1935);
    layer2_outputs(9653) <= not((layer1_outputs(5343)) or (layer1_outputs(9519)));
    layer2_outputs(9654) <= (layer1_outputs(5781)) and not (layer1_outputs(2488));
    layer2_outputs(9655) <= layer1_outputs(5495);
    layer2_outputs(9656) <= layer1_outputs(9299);
    layer2_outputs(9657) <= (layer1_outputs(3756)) and (layer1_outputs(2285));
    layer2_outputs(9658) <= layer1_outputs(6451);
    layer2_outputs(9659) <= (layer1_outputs(8781)) xor (layer1_outputs(1359));
    layer2_outputs(9660) <= '1';
    layer2_outputs(9661) <= (layer1_outputs(7413)) and (layer1_outputs(3650));
    layer2_outputs(9662) <= '1';
    layer2_outputs(9663) <= not(layer1_outputs(5653));
    layer2_outputs(9664) <= (layer1_outputs(1185)) xor (layer1_outputs(9828));
    layer2_outputs(9665) <= (layer1_outputs(7241)) and not (layer1_outputs(5044));
    layer2_outputs(9666) <= layer1_outputs(8584);
    layer2_outputs(9667) <= (layer1_outputs(6438)) xor (layer1_outputs(5551));
    layer2_outputs(9668) <= not(layer1_outputs(9223)) or (layer1_outputs(2966));
    layer2_outputs(9669) <= not((layer1_outputs(4925)) and (layer1_outputs(5463)));
    layer2_outputs(9670) <= not(layer1_outputs(6624)) or (layer1_outputs(6284));
    layer2_outputs(9671) <= layer1_outputs(8377);
    layer2_outputs(9672) <= layer1_outputs(1441);
    layer2_outputs(9673) <= (layer1_outputs(2296)) and (layer1_outputs(2362));
    layer2_outputs(9674) <= not(layer1_outputs(1113)) or (layer1_outputs(2721));
    layer2_outputs(9675) <= layer1_outputs(2927);
    layer2_outputs(9676) <= not((layer1_outputs(4947)) and (layer1_outputs(4596)));
    layer2_outputs(9677) <= (layer1_outputs(6782)) and not (layer1_outputs(5489));
    layer2_outputs(9678) <= (layer1_outputs(4925)) and not (layer1_outputs(1250));
    layer2_outputs(9679) <= not(layer1_outputs(3080));
    layer2_outputs(9680) <= not(layer1_outputs(9285)) or (layer1_outputs(4992));
    layer2_outputs(9681) <= layer1_outputs(9729);
    layer2_outputs(9682) <= not(layer1_outputs(194));
    layer2_outputs(9683) <= (layer1_outputs(4301)) xor (layer1_outputs(9400));
    layer2_outputs(9684) <= not(layer1_outputs(4692));
    layer2_outputs(9685) <= not(layer1_outputs(8491)) or (layer1_outputs(1940));
    layer2_outputs(9686) <= layer1_outputs(3857);
    layer2_outputs(9687) <= not(layer1_outputs(3273));
    layer2_outputs(9688) <= layer1_outputs(183);
    layer2_outputs(9689) <= layer1_outputs(6489);
    layer2_outputs(9690) <= not(layer1_outputs(4315)) or (layer1_outputs(2937));
    layer2_outputs(9691) <= not(layer1_outputs(8426));
    layer2_outputs(9692) <= not((layer1_outputs(7005)) and (layer1_outputs(1532)));
    layer2_outputs(9693) <= (layer1_outputs(793)) and (layer1_outputs(9561));
    layer2_outputs(9694) <= (layer1_outputs(1692)) and (layer1_outputs(2338));
    layer2_outputs(9695) <= not(layer1_outputs(3773));
    layer2_outputs(9696) <= not(layer1_outputs(6625));
    layer2_outputs(9697) <= layer1_outputs(4188);
    layer2_outputs(9698) <= not((layer1_outputs(8382)) and (layer1_outputs(509)));
    layer2_outputs(9699) <= not(layer1_outputs(6811));
    layer2_outputs(9700) <= (layer1_outputs(418)) and not (layer1_outputs(6407));
    layer2_outputs(9701) <= layer1_outputs(9694);
    layer2_outputs(9702) <= not(layer1_outputs(3259));
    layer2_outputs(9703) <= (layer1_outputs(9342)) xor (layer1_outputs(1946));
    layer2_outputs(9704) <= not((layer1_outputs(2162)) xor (layer1_outputs(6693)));
    layer2_outputs(9705) <= layer1_outputs(2520);
    layer2_outputs(9706) <= (layer1_outputs(2996)) or (layer1_outputs(2941));
    layer2_outputs(9707) <= (layer1_outputs(6269)) and (layer1_outputs(9083));
    layer2_outputs(9708) <= layer1_outputs(5847);
    layer2_outputs(9709) <= layer1_outputs(5102);
    layer2_outputs(9710) <= not(layer1_outputs(55));
    layer2_outputs(9711) <= not(layer1_outputs(4835));
    layer2_outputs(9712) <= not(layer1_outputs(7307));
    layer2_outputs(9713) <= not((layer1_outputs(750)) and (layer1_outputs(6996)));
    layer2_outputs(9714) <= (layer1_outputs(245)) and (layer1_outputs(2054));
    layer2_outputs(9715) <= not(layer1_outputs(6353)) or (layer1_outputs(9807));
    layer2_outputs(9716) <= not((layer1_outputs(3361)) xor (layer1_outputs(9858)));
    layer2_outputs(9717) <= not(layer1_outputs(7773)) or (layer1_outputs(875));
    layer2_outputs(9718) <= not(layer1_outputs(7260));
    layer2_outputs(9719) <= (layer1_outputs(8240)) xor (layer1_outputs(415));
    layer2_outputs(9720) <= (layer1_outputs(7011)) and (layer1_outputs(2081));
    layer2_outputs(9721) <= (layer1_outputs(5068)) xor (layer1_outputs(750));
    layer2_outputs(9722) <= not((layer1_outputs(6151)) or (layer1_outputs(2127)));
    layer2_outputs(9723) <= not(layer1_outputs(431)) or (layer1_outputs(5311));
    layer2_outputs(9724) <= layer1_outputs(8721);
    layer2_outputs(9725) <= not((layer1_outputs(1874)) and (layer1_outputs(5289)));
    layer2_outputs(9726) <= not(layer1_outputs(7933)) or (layer1_outputs(1655));
    layer2_outputs(9727) <= layer1_outputs(5588);
    layer2_outputs(9728) <= layer1_outputs(2339);
    layer2_outputs(9729) <= not(layer1_outputs(9821)) or (layer1_outputs(3920));
    layer2_outputs(9730) <= not(layer1_outputs(9793));
    layer2_outputs(9731) <= not(layer1_outputs(6493));
    layer2_outputs(9732) <= (layer1_outputs(3424)) and not (layer1_outputs(7201));
    layer2_outputs(9733) <= not(layer1_outputs(7817));
    layer2_outputs(9734) <= (layer1_outputs(2387)) xor (layer1_outputs(6557));
    layer2_outputs(9735) <= (layer1_outputs(4999)) xor (layer1_outputs(6090));
    layer2_outputs(9736) <= layer1_outputs(1122);
    layer2_outputs(9737) <= layer1_outputs(5577);
    layer2_outputs(9738) <= not((layer1_outputs(3173)) or (layer1_outputs(6676)));
    layer2_outputs(9739) <= not((layer1_outputs(3056)) or (layer1_outputs(9715)));
    layer2_outputs(9740) <= not((layer1_outputs(5724)) and (layer1_outputs(7917)));
    layer2_outputs(9741) <= not((layer1_outputs(5971)) or (layer1_outputs(3834)));
    layer2_outputs(9742) <= (layer1_outputs(3474)) and (layer1_outputs(2494));
    layer2_outputs(9743) <= (layer1_outputs(9956)) and not (layer1_outputs(5384));
    layer2_outputs(9744) <= not(layer1_outputs(2269));
    layer2_outputs(9745) <= not((layer1_outputs(5780)) or (layer1_outputs(3390)));
    layer2_outputs(9746) <= layer1_outputs(1239);
    layer2_outputs(9747) <= layer1_outputs(265);
    layer2_outputs(9748) <= (layer1_outputs(1687)) and not (layer1_outputs(6388));
    layer2_outputs(9749) <= not(layer1_outputs(7918));
    layer2_outputs(9750) <= (layer1_outputs(10082)) and not (layer1_outputs(6213));
    layer2_outputs(9751) <= not((layer1_outputs(9569)) and (layer1_outputs(1319)));
    layer2_outputs(9752) <= not(layer1_outputs(2847));
    layer2_outputs(9753) <= layer1_outputs(9516);
    layer2_outputs(9754) <= layer1_outputs(101);
    layer2_outputs(9755) <= layer1_outputs(5342);
    layer2_outputs(9756) <= layer1_outputs(9491);
    layer2_outputs(9757) <= not((layer1_outputs(5599)) and (layer1_outputs(2723)));
    layer2_outputs(9758) <= not(layer1_outputs(6099));
    layer2_outputs(9759) <= layer1_outputs(6897);
    layer2_outputs(9760) <= not(layer1_outputs(559));
    layer2_outputs(9761) <= layer1_outputs(6454);
    layer2_outputs(9762) <= (layer1_outputs(9389)) xor (layer1_outputs(7508));
    layer2_outputs(9763) <= not((layer1_outputs(8829)) and (layer1_outputs(6316)));
    layer2_outputs(9764) <= not(layer1_outputs(8946));
    layer2_outputs(9765) <= layer1_outputs(9437);
    layer2_outputs(9766) <= not(layer1_outputs(6253));
    layer2_outputs(9767) <= not((layer1_outputs(2606)) and (layer1_outputs(5513)));
    layer2_outputs(9768) <= not(layer1_outputs(4345));
    layer2_outputs(9769) <= not((layer1_outputs(863)) or (layer1_outputs(4773)));
    layer2_outputs(9770) <= (layer1_outputs(4600)) and not (layer1_outputs(9028));
    layer2_outputs(9771) <= layer1_outputs(5929);
    layer2_outputs(9772) <= (layer1_outputs(5554)) and (layer1_outputs(340));
    layer2_outputs(9773) <= layer1_outputs(561);
    layer2_outputs(9774) <= (layer1_outputs(3352)) and (layer1_outputs(3326));
    layer2_outputs(9775) <= not(layer1_outputs(2960));
    layer2_outputs(9776) <= not(layer1_outputs(2682));
    layer2_outputs(9777) <= layer1_outputs(1875);
    layer2_outputs(9778) <= not((layer1_outputs(4118)) or (layer1_outputs(9524)));
    layer2_outputs(9779) <= (layer1_outputs(8077)) and (layer1_outputs(10197));
    layer2_outputs(9780) <= not(layer1_outputs(5141));
    layer2_outputs(9781) <= layer1_outputs(8965);
    layer2_outputs(9782) <= not(layer1_outputs(9672));
    layer2_outputs(9783) <= layer1_outputs(6580);
    layer2_outputs(9784) <= layer1_outputs(2248);
    layer2_outputs(9785) <= layer1_outputs(1622);
    layer2_outputs(9786) <= not(layer1_outputs(7708)) or (layer1_outputs(7949));
    layer2_outputs(9787) <= not((layer1_outputs(6213)) and (layer1_outputs(2400)));
    layer2_outputs(9788) <= (layer1_outputs(6782)) xor (layer1_outputs(563));
    layer2_outputs(9789) <= layer1_outputs(3586);
    layer2_outputs(9790) <= layer1_outputs(3697);
    layer2_outputs(9791) <= (layer1_outputs(5942)) xor (layer1_outputs(1002));
    layer2_outputs(9792) <= (layer1_outputs(5857)) and not (layer1_outputs(37));
    layer2_outputs(9793) <= layer1_outputs(3305);
    layer2_outputs(9794) <= not(layer1_outputs(7269));
    layer2_outputs(9795) <= (layer1_outputs(3024)) or (layer1_outputs(529));
    layer2_outputs(9796) <= layer1_outputs(4666);
    layer2_outputs(9797) <= not(layer1_outputs(9831));
    layer2_outputs(9798) <= layer1_outputs(7471);
    layer2_outputs(9799) <= layer1_outputs(4318);
    layer2_outputs(9800) <= (layer1_outputs(2601)) xor (layer1_outputs(1854));
    layer2_outputs(9801) <= layer1_outputs(1036);
    layer2_outputs(9802) <= not(layer1_outputs(3291)) or (layer1_outputs(6609));
    layer2_outputs(9803) <= layer1_outputs(10026);
    layer2_outputs(9804) <= not(layer1_outputs(8608));
    layer2_outputs(9805) <= not(layer1_outputs(1884)) or (layer1_outputs(7193));
    layer2_outputs(9806) <= not(layer1_outputs(1604));
    layer2_outputs(9807) <= not((layer1_outputs(7973)) xor (layer1_outputs(3786)));
    layer2_outputs(9808) <= layer1_outputs(5104);
    layer2_outputs(9809) <= not(layer1_outputs(6399));
    layer2_outputs(9810) <= not(layer1_outputs(8279));
    layer2_outputs(9811) <= not(layer1_outputs(2982)) or (layer1_outputs(4705));
    layer2_outputs(9812) <= not(layer1_outputs(4830));
    layer2_outputs(9813) <= not(layer1_outputs(9942));
    layer2_outputs(9814) <= (layer1_outputs(9032)) and (layer1_outputs(1065));
    layer2_outputs(9815) <= layer1_outputs(2858);
    layer2_outputs(9816) <= (layer1_outputs(6788)) and not (layer1_outputs(865));
    layer2_outputs(9817) <= (layer1_outputs(3978)) and not (layer1_outputs(4927));
    layer2_outputs(9818) <= not(layer1_outputs(791));
    layer2_outputs(9819) <= not(layer1_outputs(9860));
    layer2_outputs(9820) <= (layer1_outputs(1871)) and (layer1_outputs(8394));
    layer2_outputs(9821) <= not(layer1_outputs(2425));
    layer2_outputs(9822) <= not((layer1_outputs(5685)) or (layer1_outputs(6416)));
    layer2_outputs(9823) <= not(layer1_outputs(907));
    layer2_outputs(9824) <= not((layer1_outputs(794)) and (layer1_outputs(8382)));
    layer2_outputs(9825) <= (layer1_outputs(19)) or (layer1_outputs(6691));
    layer2_outputs(9826) <= (layer1_outputs(1156)) xor (layer1_outputs(6503));
    layer2_outputs(9827) <= (layer1_outputs(7324)) and (layer1_outputs(4292));
    layer2_outputs(9828) <= layer1_outputs(8172);
    layer2_outputs(9829) <= not(layer1_outputs(8120));
    layer2_outputs(9830) <= not(layer1_outputs(7634));
    layer2_outputs(9831) <= (layer1_outputs(267)) xor (layer1_outputs(3554));
    layer2_outputs(9832) <= layer1_outputs(3781);
    layer2_outputs(9833) <= not((layer1_outputs(10148)) xor (layer1_outputs(80)));
    layer2_outputs(9834) <= not(layer1_outputs(9913));
    layer2_outputs(9835) <= layer1_outputs(9171);
    layer2_outputs(9836) <= not((layer1_outputs(3482)) xor (layer1_outputs(4755)));
    layer2_outputs(9837) <= not(layer1_outputs(6049));
    layer2_outputs(9838) <= layer1_outputs(5897);
    layer2_outputs(9839) <= not(layer1_outputs(5862));
    layer2_outputs(9840) <= (layer1_outputs(4218)) and not (layer1_outputs(7807));
    layer2_outputs(9841) <= not((layer1_outputs(772)) xor (layer1_outputs(8226)));
    layer2_outputs(9842) <= (layer1_outputs(8242)) and not (layer1_outputs(946));
    layer2_outputs(9843) <= not(layer1_outputs(2239)) or (layer1_outputs(9569));
    layer2_outputs(9844) <= layer1_outputs(7748);
    layer2_outputs(9845) <= layer1_outputs(9619);
    layer2_outputs(9846) <= layer1_outputs(4669);
    layer2_outputs(9847) <= not((layer1_outputs(7593)) or (layer1_outputs(6300)));
    layer2_outputs(9848) <= not(layer1_outputs(2200));
    layer2_outputs(9849) <= not(layer1_outputs(9306));
    layer2_outputs(9850) <= not(layer1_outputs(1433));
    layer2_outputs(9851) <= layer1_outputs(8358);
    layer2_outputs(9852) <= not(layer1_outputs(10080));
    layer2_outputs(9853) <= layer1_outputs(7663);
    layer2_outputs(9854) <= not((layer1_outputs(7835)) and (layer1_outputs(3909)));
    layer2_outputs(9855) <= not(layer1_outputs(9729));
    layer2_outputs(9856) <= not(layer1_outputs(1025));
    layer2_outputs(9857) <= not(layer1_outputs(5925));
    layer2_outputs(9858) <= not(layer1_outputs(8379));
    layer2_outputs(9859) <= not((layer1_outputs(5179)) xor (layer1_outputs(2404)));
    layer2_outputs(9860) <= (layer1_outputs(5070)) and (layer1_outputs(9448));
    layer2_outputs(9861) <= not(layer1_outputs(6097));
    layer2_outputs(9862) <= not((layer1_outputs(930)) and (layer1_outputs(5432)));
    layer2_outputs(9863) <= not(layer1_outputs(281));
    layer2_outputs(9864) <= not(layer1_outputs(1744)) or (layer1_outputs(4523));
    layer2_outputs(9865) <= (layer1_outputs(8533)) and not (layer1_outputs(6135));
    layer2_outputs(9866) <= not((layer1_outputs(8040)) xor (layer1_outputs(7434)));
    layer2_outputs(9867) <= layer1_outputs(2206);
    layer2_outputs(9868) <= (layer1_outputs(3645)) and (layer1_outputs(4013));
    layer2_outputs(9869) <= layer1_outputs(1624);
    layer2_outputs(9870) <= not((layer1_outputs(227)) xor (layer1_outputs(8609)));
    layer2_outputs(9871) <= not(layer1_outputs(7924)) or (layer1_outputs(6744));
    layer2_outputs(9872) <= (layer1_outputs(9182)) xor (layer1_outputs(7385));
    layer2_outputs(9873) <= not(layer1_outputs(1128));
    layer2_outputs(9874) <= not(layer1_outputs(3937));
    layer2_outputs(9875) <= layer1_outputs(3326);
    layer2_outputs(9876) <= layer1_outputs(890);
    layer2_outputs(9877) <= layer1_outputs(3812);
    layer2_outputs(9878) <= not(layer1_outputs(334)) or (layer1_outputs(1977));
    layer2_outputs(9879) <= (layer1_outputs(2679)) and (layer1_outputs(2444));
    layer2_outputs(9880) <= not((layer1_outputs(1027)) and (layer1_outputs(9871)));
    layer2_outputs(9881) <= not(layer1_outputs(5928)) or (layer1_outputs(8694));
    layer2_outputs(9882) <= layer1_outputs(1569);
    layer2_outputs(9883) <= not(layer1_outputs(4778));
    layer2_outputs(9884) <= '0';
    layer2_outputs(9885) <= layer1_outputs(8971);
    layer2_outputs(9886) <= layer1_outputs(8430);
    layer2_outputs(9887) <= not(layer1_outputs(4344));
    layer2_outputs(9888) <= not(layer1_outputs(1223)) or (layer1_outputs(1277));
    layer2_outputs(9889) <= not(layer1_outputs(2940));
    layer2_outputs(9890) <= (layer1_outputs(4713)) and (layer1_outputs(1152));
    layer2_outputs(9891) <= (layer1_outputs(8508)) and (layer1_outputs(7379));
    layer2_outputs(9892) <= not((layer1_outputs(24)) and (layer1_outputs(8486)));
    layer2_outputs(9893) <= not(layer1_outputs(9025)) or (layer1_outputs(1147));
    layer2_outputs(9894) <= not(layer1_outputs(1845));
    layer2_outputs(9895) <= not(layer1_outputs(3448)) or (layer1_outputs(6917));
    layer2_outputs(9896) <= not(layer1_outputs(5832));
    layer2_outputs(9897) <= not(layer1_outputs(6740));
    layer2_outputs(9898) <= not(layer1_outputs(8390));
    layer2_outputs(9899) <= not((layer1_outputs(4906)) or (layer1_outputs(7554)));
    layer2_outputs(9900) <= (layer1_outputs(1320)) and not (layer1_outputs(134));
    layer2_outputs(9901) <= not((layer1_outputs(8766)) and (layer1_outputs(1843)));
    layer2_outputs(9902) <= not(layer1_outputs(6034));
    layer2_outputs(9903) <= not((layer1_outputs(7668)) xor (layer1_outputs(10218)));
    layer2_outputs(9904) <= (layer1_outputs(6475)) and not (layer1_outputs(6122));
    layer2_outputs(9905) <= not(layer1_outputs(9591)) or (layer1_outputs(3040));
    layer2_outputs(9906) <= not(layer1_outputs(1670));
    layer2_outputs(9907) <= (layer1_outputs(6614)) xor (layer1_outputs(3742));
    layer2_outputs(9908) <= not(layer1_outputs(3830));
    layer2_outputs(9909) <= not(layer1_outputs(3957)) or (layer1_outputs(4933));
    layer2_outputs(9910) <= layer1_outputs(661);
    layer2_outputs(9911) <= layer1_outputs(456);
    layer2_outputs(9912) <= layer1_outputs(9935);
    layer2_outputs(9913) <= not((layer1_outputs(5089)) and (layer1_outputs(9632)));
    layer2_outputs(9914) <= not(layer1_outputs(299));
    layer2_outputs(9915) <= '0';
    layer2_outputs(9916) <= (layer1_outputs(2379)) and not (layer1_outputs(3451));
    layer2_outputs(9917) <= (layer1_outputs(1950)) and not (layer1_outputs(8548));
    layer2_outputs(9918) <= not(layer1_outputs(9342));
    layer2_outputs(9919) <= not(layer1_outputs(4162));
    layer2_outputs(9920) <= not(layer1_outputs(3048)) or (layer1_outputs(7350));
    layer2_outputs(9921) <= not(layer1_outputs(3897)) or (layer1_outputs(7085));
    layer2_outputs(9922) <= not(layer1_outputs(9222));
    layer2_outputs(9923) <= not(layer1_outputs(6321));
    layer2_outputs(9924) <= layer1_outputs(1456);
    layer2_outputs(9925) <= not(layer1_outputs(2768));
    layer2_outputs(9926) <= (layer1_outputs(1474)) xor (layer1_outputs(1119));
    layer2_outputs(9927) <= (layer1_outputs(8091)) and (layer1_outputs(380));
    layer2_outputs(9928) <= (layer1_outputs(9933)) or (layer1_outputs(4542));
    layer2_outputs(9929) <= not(layer1_outputs(1841)) or (layer1_outputs(2711));
    layer2_outputs(9930) <= (layer1_outputs(7760)) xor (layer1_outputs(1522));
    layer2_outputs(9931) <= (layer1_outputs(89)) or (layer1_outputs(10211));
    layer2_outputs(9932) <= not(layer1_outputs(774));
    layer2_outputs(9933) <= not(layer1_outputs(10157)) or (layer1_outputs(7363));
    layer2_outputs(9934) <= not((layer1_outputs(1602)) or (layer1_outputs(6016)));
    layer2_outputs(9935) <= '0';
    layer2_outputs(9936) <= not((layer1_outputs(4160)) or (layer1_outputs(1711)));
    layer2_outputs(9937) <= not(layer1_outputs(2920));
    layer2_outputs(9938) <= (layer1_outputs(1787)) or (layer1_outputs(3561));
    layer2_outputs(9939) <= (layer1_outputs(5941)) xor (layer1_outputs(2757));
    layer2_outputs(9940) <= (layer1_outputs(6161)) xor (layer1_outputs(2155));
    layer2_outputs(9941) <= not(layer1_outputs(4646));
    layer2_outputs(9942) <= layer1_outputs(2498);
    layer2_outputs(9943) <= not(layer1_outputs(4820)) or (layer1_outputs(9868));
    layer2_outputs(9944) <= layer1_outputs(5387);
    layer2_outputs(9945) <= layer1_outputs(143);
    layer2_outputs(9946) <= layer1_outputs(1915);
    layer2_outputs(9947) <= not(layer1_outputs(9949));
    layer2_outputs(9948) <= layer1_outputs(535);
    layer2_outputs(9949) <= (layer1_outputs(403)) and not (layer1_outputs(3222));
    layer2_outputs(9950) <= (layer1_outputs(4210)) xor (layer1_outputs(7980));
    layer2_outputs(9951) <= not((layer1_outputs(6824)) xor (layer1_outputs(171)));
    layer2_outputs(9952) <= layer1_outputs(9292);
    layer2_outputs(9953) <= not(layer1_outputs(7079));
    layer2_outputs(9954) <= (layer1_outputs(4514)) and not (layer1_outputs(4909));
    layer2_outputs(9955) <= (layer1_outputs(4061)) xor (layer1_outputs(8489));
    layer2_outputs(9956) <= not((layer1_outputs(481)) xor (layer1_outputs(398)));
    layer2_outputs(9957) <= (layer1_outputs(6854)) or (layer1_outputs(8280));
    layer2_outputs(9958) <= layer1_outputs(7251);
    layer2_outputs(9959) <= not(layer1_outputs(4308)) or (layer1_outputs(7210));
    layer2_outputs(9960) <= not(layer1_outputs(8324)) or (layer1_outputs(8856));
    layer2_outputs(9961) <= layer1_outputs(9189);
    layer2_outputs(9962) <= not(layer1_outputs(9585));
    layer2_outputs(9963) <= '0';
    layer2_outputs(9964) <= not((layer1_outputs(1916)) xor (layer1_outputs(1484)));
    layer2_outputs(9965) <= not(layer1_outputs(2179)) or (layer1_outputs(5610));
    layer2_outputs(9966) <= layer1_outputs(2844);
    layer2_outputs(9967) <= not((layer1_outputs(1944)) xor (layer1_outputs(5573)));
    layer2_outputs(9968) <= (layer1_outputs(7635)) and not (layer1_outputs(9487));
    layer2_outputs(9969) <= layer1_outputs(5418);
    layer2_outputs(9970) <= not(layer1_outputs(4686));
    layer2_outputs(9971) <= layer1_outputs(9604);
    layer2_outputs(9972) <= not(layer1_outputs(2311)) or (layer1_outputs(3085));
    layer2_outputs(9973) <= not(layer1_outputs(1218));
    layer2_outputs(9974) <= layer1_outputs(1807);
    layer2_outputs(9975) <= (layer1_outputs(3133)) or (layer1_outputs(1787));
    layer2_outputs(9976) <= not(layer1_outputs(8505));
    layer2_outputs(9977) <= not(layer1_outputs(4435));
    layer2_outputs(9978) <= (layer1_outputs(9275)) or (layer1_outputs(3966));
    layer2_outputs(9979) <= (layer1_outputs(1322)) and not (layer1_outputs(6182));
    layer2_outputs(9980) <= not(layer1_outputs(5686)) or (layer1_outputs(8058));
    layer2_outputs(9981) <= layer1_outputs(3250);
    layer2_outputs(9982) <= not(layer1_outputs(1194));
    layer2_outputs(9983) <= (layer1_outputs(6849)) xor (layer1_outputs(9247));
    layer2_outputs(9984) <= not(layer1_outputs(3719));
    layer2_outputs(9985) <= not((layer1_outputs(4704)) or (layer1_outputs(5484)));
    layer2_outputs(9986) <= layer1_outputs(6379);
    layer2_outputs(9987) <= (layer1_outputs(4355)) and (layer1_outputs(1465));
    layer2_outputs(9988) <= (layer1_outputs(7245)) and (layer1_outputs(7091));
    layer2_outputs(9989) <= not((layer1_outputs(4370)) xor (layer1_outputs(2612)));
    layer2_outputs(9990) <= (layer1_outputs(8645)) and not (layer1_outputs(6965));
    layer2_outputs(9991) <= not(layer1_outputs(9399));
    layer2_outputs(9992) <= (layer1_outputs(9919)) xor (layer1_outputs(654));
    layer2_outputs(9993) <= not(layer1_outputs(6308));
    layer2_outputs(9994) <= layer1_outputs(4867);
    layer2_outputs(9995) <= not(layer1_outputs(2872)) or (layer1_outputs(438));
    layer2_outputs(9996) <= not(layer1_outputs(7022));
    layer2_outputs(9997) <= layer1_outputs(5236);
    layer2_outputs(9998) <= (layer1_outputs(5059)) and not (layer1_outputs(1002));
    layer2_outputs(9999) <= (layer1_outputs(3197)) and not (layer1_outputs(1533));
    layer2_outputs(10000) <= (layer1_outputs(5487)) and not (layer1_outputs(5957));
    layer2_outputs(10001) <= not((layer1_outputs(1093)) or (layer1_outputs(1008)));
    layer2_outputs(10002) <= not((layer1_outputs(6186)) or (layer1_outputs(4066)));
    layer2_outputs(10003) <= not((layer1_outputs(6005)) or (layer1_outputs(7580)));
    layer2_outputs(10004) <= not(layer1_outputs(5774));
    layer2_outputs(10005) <= layer1_outputs(7430);
    layer2_outputs(10006) <= not(layer1_outputs(1447));
    layer2_outputs(10007) <= layer1_outputs(4764);
    layer2_outputs(10008) <= not((layer1_outputs(439)) or (layer1_outputs(5391)));
    layer2_outputs(10009) <= not(layer1_outputs(6541));
    layer2_outputs(10010) <= not(layer1_outputs(7794));
    layer2_outputs(10011) <= layer1_outputs(5658);
    layer2_outputs(10012) <= layer1_outputs(7890);
    layer2_outputs(10013) <= '0';
    layer2_outputs(10014) <= '1';
    layer2_outputs(10015) <= layer1_outputs(454);
    layer2_outputs(10016) <= not((layer1_outputs(3299)) xor (layer1_outputs(2390)));
    layer2_outputs(10017) <= layer1_outputs(3691);
    layer2_outputs(10018) <= not(layer1_outputs(2913)) or (layer1_outputs(8848));
    layer2_outputs(10019) <= layer1_outputs(8830);
    layer2_outputs(10020) <= (layer1_outputs(765)) and not (layer1_outputs(5841));
    layer2_outputs(10021) <= layer1_outputs(7494);
    layer2_outputs(10022) <= not((layer1_outputs(263)) or (layer1_outputs(7369)));
    layer2_outputs(10023) <= not((layer1_outputs(4471)) xor (layer1_outputs(3616)));
    layer2_outputs(10024) <= not(layer1_outputs(8805)) or (layer1_outputs(5115));
    layer2_outputs(10025) <= (layer1_outputs(6830)) xor (layer1_outputs(9080));
    layer2_outputs(10026) <= not((layer1_outputs(2408)) and (layer1_outputs(727)));
    layer2_outputs(10027) <= not(layer1_outputs(6168));
    layer2_outputs(10028) <= (layer1_outputs(8187)) and (layer1_outputs(8786));
    layer2_outputs(10029) <= not((layer1_outputs(1299)) and (layer1_outputs(7164)));
    layer2_outputs(10030) <= layer1_outputs(1210);
    layer2_outputs(10031) <= (layer1_outputs(4113)) or (layer1_outputs(1417));
    layer2_outputs(10032) <= not(layer1_outputs(5065));
    layer2_outputs(10033) <= not((layer1_outputs(2200)) or (layer1_outputs(3873)));
    layer2_outputs(10034) <= not(layer1_outputs(7120));
    layer2_outputs(10035) <= not(layer1_outputs(9283));
    layer2_outputs(10036) <= (layer1_outputs(8239)) and not (layer1_outputs(8808));
    layer2_outputs(10037) <= not(layer1_outputs(2942)) or (layer1_outputs(7334));
    layer2_outputs(10038) <= layer1_outputs(3565);
    layer2_outputs(10039) <= layer1_outputs(137);
    layer2_outputs(10040) <= not(layer1_outputs(334));
    layer2_outputs(10041) <= layer1_outputs(3529);
    layer2_outputs(10042) <= (layer1_outputs(7770)) or (layer1_outputs(9883));
    layer2_outputs(10043) <= layer1_outputs(9613);
    layer2_outputs(10044) <= not(layer1_outputs(2173));
    layer2_outputs(10045) <= not((layer1_outputs(7373)) xor (layer1_outputs(54)));
    layer2_outputs(10046) <= not(layer1_outputs(8210));
    layer2_outputs(10047) <= layer1_outputs(3143);
    layer2_outputs(10048) <= (layer1_outputs(1092)) and not (layer1_outputs(1415));
    layer2_outputs(10049) <= not(layer1_outputs(6867));
    layer2_outputs(10050) <= layer1_outputs(8822);
    layer2_outputs(10051) <= (layer1_outputs(174)) and not (layer1_outputs(7263));
    layer2_outputs(10052) <= not(layer1_outputs(8373));
    layer2_outputs(10053) <= (layer1_outputs(896)) or (layer1_outputs(31));
    layer2_outputs(10054) <= (layer1_outputs(600)) and not (layer1_outputs(8552));
    layer2_outputs(10055) <= (layer1_outputs(9493)) and (layer1_outputs(9368));
    layer2_outputs(10056) <= not((layer1_outputs(4022)) or (layer1_outputs(3851)));
    layer2_outputs(10057) <= (layer1_outputs(4091)) and (layer1_outputs(4411));
    layer2_outputs(10058) <= layer1_outputs(2578);
    layer2_outputs(10059) <= not(layer1_outputs(8168)) or (layer1_outputs(10235));
    layer2_outputs(10060) <= (layer1_outputs(6225)) or (layer1_outputs(5079));
    layer2_outputs(10061) <= not(layer1_outputs(9266));
    layer2_outputs(10062) <= not((layer1_outputs(3465)) and (layer1_outputs(4432)));
    layer2_outputs(10063) <= not(layer1_outputs(729)) or (layer1_outputs(7278));
    layer2_outputs(10064) <= layer1_outputs(9362);
    layer2_outputs(10065) <= not(layer1_outputs(4662));
    layer2_outputs(10066) <= (layer1_outputs(8103)) and not (layer1_outputs(7247));
    layer2_outputs(10067) <= layer1_outputs(3053);
    layer2_outputs(10068) <= layer1_outputs(6992);
    layer2_outputs(10069) <= layer1_outputs(7412);
    layer2_outputs(10070) <= not(layer1_outputs(1115));
    layer2_outputs(10071) <= not(layer1_outputs(5004));
    layer2_outputs(10072) <= layer1_outputs(1564);
    layer2_outputs(10073) <= (layer1_outputs(1524)) and not (layer1_outputs(3706));
    layer2_outputs(10074) <= not((layer1_outputs(3110)) xor (layer1_outputs(8626)));
    layer2_outputs(10075) <= not(layer1_outputs(6054));
    layer2_outputs(10076) <= layer1_outputs(7495);
    layer2_outputs(10077) <= (layer1_outputs(9965)) or (layer1_outputs(9982));
    layer2_outputs(10078) <= not(layer1_outputs(544));
    layer2_outputs(10079) <= (layer1_outputs(8144)) xor (layer1_outputs(9556));
    layer2_outputs(10080) <= not((layer1_outputs(7553)) xor (layer1_outputs(4866)));
    layer2_outputs(10081) <= '0';
    layer2_outputs(10082) <= not((layer1_outputs(9461)) xor (layer1_outputs(2249)));
    layer2_outputs(10083) <= not((layer1_outputs(7147)) or (layer1_outputs(3968)));
    layer2_outputs(10084) <= layer1_outputs(5698);
    layer2_outputs(10085) <= (layer1_outputs(4112)) xor (layer1_outputs(10039));
    layer2_outputs(10086) <= (layer1_outputs(9747)) and not (layer1_outputs(9889));
    layer2_outputs(10087) <= (layer1_outputs(8606)) and not (layer1_outputs(3299));
    layer2_outputs(10088) <= (layer1_outputs(3789)) and not (layer1_outputs(6924));
    layer2_outputs(10089) <= not(layer1_outputs(2767)) or (layer1_outputs(4387));
    layer2_outputs(10090) <= layer1_outputs(8908);
    layer2_outputs(10091) <= (layer1_outputs(6711)) and not (layer1_outputs(8262));
    layer2_outputs(10092) <= not(layer1_outputs(6688));
    layer2_outputs(10093) <= not(layer1_outputs(251)) or (layer1_outputs(9906));
    layer2_outputs(10094) <= not((layer1_outputs(965)) or (layer1_outputs(3503)));
    layer2_outputs(10095) <= layer1_outputs(8742);
    layer2_outputs(10096) <= not((layer1_outputs(6227)) xor (layer1_outputs(3958)));
    layer2_outputs(10097) <= (layer1_outputs(4395)) and (layer1_outputs(6948));
    layer2_outputs(10098) <= not(layer1_outputs(8447));
    layer2_outputs(10099) <= layer1_outputs(4817);
    layer2_outputs(10100) <= layer1_outputs(9468);
    layer2_outputs(10101) <= not(layer1_outputs(6726));
    layer2_outputs(10102) <= (layer1_outputs(6926)) and (layer1_outputs(8404));
    layer2_outputs(10103) <= layer1_outputs(40);
    layer2_outputs(10104) <= layer1_outputs(5230);
    layer2_outputs(10105) <= layer1_outputs(6769);
    layer2_outputs(10106) <= layer1_outputs(9291);
    layer2_outputs(10107) <= not(layer1_outputs(8099));
    layer2_outputs(10108) <= not(layer1_outputs(5874));
    layer2_outputs(10109) <= (layer1_outputs(9874)) xor (layer1_outputs(2120));
    layer2_outputs(10110) <= layer1_outputs(2858);
    layer2_outputs(10111) <= not(layer1_outputs(6153));
    layer2_outputs(10112) <= not(layer1_outputs(3732)) or (layer1_outputs(5272));
    layer2_outputs(10113) <= (layer1_outputs(8086)) or (layer1_outputs(1955));
    layer2_outputs(10114) <= not(layer1_outputs(7485)) or (layer1_outputs(7986));
    layer2_outputs(10115) <= (layer1_outputs(6292)) and (layer1_outputs(10215));
    layer2_outputs(10116) <= (layer1_outputs(7560)) xor (layer1_outputs(9306));
    layer2_outputs(10117) <= (layer1_outputs(4812)) and not (layer1_outputs(5033));
    layer2_outputs(10118) <= (layer1_outputs(8570)) xor (layer1_outputs(2429));
    layer2_outputs(10119) <= not(layer1_outputs(2624)) or (layer1_outputs(9436));
    layer2_outputs(10120) <= layer1_outputs(9499);
    layer2_outputs(10121) <= '0';
    layer2_outputs(10122) <= not(layer1_outputs(8078));
    layer2_outputs(10123) <= (layer1_outputs(3058)) and not (layer1_outputs(9772));
    layer2_outputs(10124) <= layer1_outputs(5313);
    layer2_outputs(10125) <= (layer1_outputs(6750)) or (layer1_outputs(5853));
    layer2_outputs(10126) <= not(layer1_outputs(4643));
    layer2_outputs(10127) <= not(layer1_outputs(4896));
    layer2_outputs(10128) <= not((layer1_outputs(132)) and (layer1_outputs(4757)));
    layer2_outputs(10129) <= not(layer1_outputs(9756));
    layer2_outputs(10130) <= not((layer1_outputs(3872)) and (layer1_outputs(1205)));
    layer2_outputs(10131) <= not(layer1_outputs(9531));
    layer2_outputs(10132) <= not(layer1_outputs(2993));
    layer2_outputs(10133) <= layer1_outputs(394);
    layer2_outputs(10134) <= not((layer1_outputs(7968)) or (layer1_outputs(7313)));
    layer2_outputs(10135) <= (layer1_outputs(9377)) xor (layer1_outputs(1975));
    layer2_outputs(10136) <= not(layer1_outputs(8765));
    layer2_outputs(10137) <= not((layer1_outputs(8073)) and (layer1_outputs(7840)));
    layer2_outputs(10138) <= (layer1_outputs(1376)) and not (layer1_outputs(8187));
    layer2_outputs(10139) <= not(layer1_outputs(2586)) or (layer1_outputs(7311));
    layer2_outputs(10140) <= '1';
    layer2_outputs(10141) <= (layer1_outputs(5567)) and not (layer1_outputs(1916));
    layer2_outputs(10142) <= not(layer1_outputs(8737));
    layer2_outputs(10143) <= not(layer1_outputs(2855)) or (layer1_outputs(1577));
    layer2_outputs(10144) <= not((layer1_outputs(2245)) and (layer1_outputs(8444)));
    layer2_outputs(10145) <= not(layer1_outputs(3273));
    layer2_outputs(10146) <= not(layer1_outputs(8904));
    layer2_outputs(10147) <= (layer1_outputs(4476)) and not (layer1_outputs(2015));
    layer2_outputs(10148) <= layer1_outputs(2613);
    layer2_outputs(10149) <= not(layer1_outputs(7671));
    layer2_outputs(10150) <= not(layer1_outputs(955));
    layer2_outputs(10151) <= (layer1_outputs(2970)) and not (layer1_outputs(914));
    layer2_outputs(10152) <= not(layer1_outputs(8418));
    layer2_outputs(10153) <= (layer1_outputs(3695)) xor (layer1_outputs(2213));
    layer2_outputs(10154) <= (layer1_outputs(9295)) xor (layer1_outputs(3981));
    layer2_outputs(10155) <= layer1_outputs(3643);
    layer2_outputs(10156) <= not((layer1_outputs(7642)) xor (layer1_outputs(7900)));
    layer2_outputs(10157) <= layer1_outputs(8371);
    layer2_outputs(10158) <= not((layer1_outputs(547)) xor (layer1_outputs(8707)));
    layer2_outputs(10159) <= not(layer1_outputs(7532)) or (layer1_outputs(5495));
    layer2_outputs(10160) <= not((layer1_outputs(5419)) and (layer1_outputs(4360)));
    layer2_outputs(10161) <= not((layer1_outputs(8581)) or (layer1_outputs(5204)));
    layer2_outputs(10162) <= not(layer1_outputs(6053)) or (layer1_outputs(8376));
    layer2_outputs(10163) <= layer1_outputs(4729);
    layer2_outputs(10164) <= (layer1_outputs(3372)) and not (layer1_outputs(5200));
    layer2_outputs(10165) <= not((layer1_outputs(3008)) and (layer1_outputs(8626)));
    layer2_outputs(10166) <= (layer1_outputs(2250)) and not (layer1_outputs(8847));
    layer2_outputs(10167) <= not(layer1_outputs(2539));
    layer2_outputs(10168) <= (layer1_outputs(6609)) and not (layer1_outputs(111));
    layer2_outputs(10169) <= not((layer1_outputs(5939)) and (layer1_outputs(9733)));
    layer2_outputs(10170) <= not(layer1_outputs(2542)) or (layer1_outputs(2519));
    layer2_outputs(10171) <= not(layer1_outputs(4069));
    layer2_outputs(10172) <= '0';
    layer2_outputs(10173) <= (layer1_outputs(4356)) xor (layer1_outputs(2467));
    layer2_outputs(10174) <= layer1_outputs(2976);
    layer2_outputs(10175) <= not((layer1_outputs(4083)) xor (layer1_outputs(9129)));
    layer2_outputs(10176) <= not(layer1_outputs(3986));
    layer2_outputs(10177) <= (layer1_outputs(9262)) and (layer1_outputs(8972));
    layer2_outputs(10178) <= not(layer1_outputs(5853));
    layer2_outputs(10179) <= layer1_outputs(1045);
    layer2_outputs(10180) <= not(layer1_outputs(9514)) or (layer1_outputs(2800));
    layer2_outputs(10181) <= (layer1_outputs(5822)) xor (layer1_outputs(411));
    layer2_outputs(10182) <= layer1_outputs(2011);
    layer2_outputs(10183) <= not(layer1_outputs(3453)) or (layer1_outputs(5761));
    layer2_outputs(10184) <= not((layer1_outputs(1018)) and (layer1_outputs(9518)));
    layer2_outputs(10185) <= not((layer1_outputs(2158)) xor (layer1_outputs(3647)));
    layer2_outputs(10186) <= not(layer1_outputs(10078));
    layer2_outputs(10187) <= layer1_outputs(3696);
    layer2_outputs(10188) <= (layer1_outputs(10037)) xor (layer1_outputs(4840));
    layer2_outputs(10189) <= not(layer1_outputs(5226));
    layer2_outputs(10190) <= (layer1_outputs(258)) and not (layer1_outputs(3149));
    layer2_outputs(10191) <= not((layer1_outputs(9148)) xor (layer1_outputs(8597)));
    layer2_outputs(10192) <= layer1_outputs(9043);
    layer2_outputs(10193) <= (layer1_outputs(2312)) and not (layer1_outputs(8646));
    layer2_outputs(10194) <= not(layer1_outputs(5097));
    layer2_outputs(10195) <= (layer1_outputs(1215)) or (layer1_outputs(8817));
    layer2_outputs(10196) <= not((layer1_outputs(6629)) xor (layer1_outputs(6098)));
    layer2_outputs(10197) <= (layer1_outputs(422)) and not (layer1_outputs(3719));
    layer2_outputs(10198) <= not((layer1_outputs(1306)) xor (layer1_outputs(7387)));
    layer2_outputs(10199) <= (layer1_outputs(407)) or (layer1_outputs(6835));
    layer2_outputs(10200) <= not(layer1_outputs(8699)) or (layer1_outputs(4135));
    layer2_outputs(10201) <= not((layer1_outputs(6573)) or (layer1_outputs(657)));
    layer2_outputs(10202) <= layer1_outputs(5655);
    layer2_outputs(10203) <= layer1_outputs(3285);
    layer2_outputs(10204) <= not((layer1_outputs(7977)) and (layer1_outputs(9157)));
    layer2_outputs(10205) <= not(layer1_outputs(4821)) or (layer1_outputs(6130));
    layer2_outputs(10206) <= not(layer1_outputs(3578));
    layer2_outputs(10207) <= not((layer1_outputs(4539)) and (layer1_outputs(6492)));
    layer2_outputs(10208) <= layer1_outputs(4269);
    layer2_outputs(10209) <= not(layer1_outputs(2845));
    layer2_outputs(10210) <= not((layer1_outputs(6711)) and (layer1_outputs(8345)));
    layer2_outputs(10211) <= not((layer1_outputs(6839)) xor (layer1_outputs(589)));
    layer2_outputs(10212) <= not(layer1_outputs(9369)) or (layer1_outputs(2358));
    layer2_outputs(10213) <= not(layer1_outputs(2046));
    layer2_outputs(10214) <= (layer1_outputs(2350)) and not (layer1_outputs(4990));
    layer2_outputs(10215) <= layer1_outputs(9029);
    layer2_outputs(10216) <= layer1_outputs(6146);
    layer2_outputs(10217) <= (layer1_outputs(1685)) and not (layer1_outputs(3914));
    layer2_outputs(10218) <= layer1_outputs(2716);
    layer2_outputs(10219) <= not((layer1_outputs(3999)) xor (layer1_outputs(6111)));
    layer2_outputs(10220) <= not((layer1_outputs(4323)) or (layer1_outputs(2840)));
    layer2_outputs(10221) <= not((layer1_outputs(1759)) xor (layer1_outputs(3495)));
    layer2_outputs(10222) <= (layer1_outputs(7540)) and not (layer1_outputs(9472));
    layer2_outputs(10223) <= '1';
    layer2_outputs(10224) <= layer1_outputs(1379);
    layer2_outputs(10225) <= not(layer1_outputs(3433));
    layer2_outputs(10226) <= (layer1_outputs(6382)) and not (layer1_outputs(2673));
    layer2_outputs(10227) <= layer1_outputs(9513);
    layer2_outputs(10228) <= (layer1_outputs(2256)) and not (layer1_outputs(4319));
    layer2_outputs(10229) <= not((layer1_outputs(3232)) or (layer1_outputs(3146)));
    layer2_outputs(10230) <= (layer1_outputs(3497)) and not (layer1_outputs(5746));
    layer2_outputs(10231) <= not(layer1_outputs(8815)) or (layer1_outputs(3858));
    layer2_outputs(10232) <= not(layer1_outputs(5887));
    layer2_outputs(10233) <= (layer1_outputs(7820)) and not (layer1_outputs(5400));
    layer2_outputs(10234) <= layer1_outputs(1479);
    layer2_outputs(10235) <= (layer1_outputs(4039)) xor (layer1_outputs(7711));
    layer2_outputs(10236) <= not(layer1_outputs(5734));
    layer2_outputs(10237) <= not(layer1_outputs(5710)) or (layer1_outputs(4990));
    layer2_outputs(10238) <= not(layer1_outputs(6263)) or (layer1_outputs(2399));
    layer2_outputs(10239) <= not(layer1_outputs(4971)) or (layer1_outputs(4400));
    outputs(0) <= not(layer2_outputs(2099));
    outputs(1) <= layer2_outputs(723);
    outputs(2) <= layer2_outputs(2390);
    outputs(3) <= not((layer2_outputs(9594)) and (layer2_outputs(3751)));
    outputs(4) <= layer2_outputs(1428);
    outputs(5) <= (layer2_outputs(7725)) and (layer2_outputs(1846));
    outputs(6) <= (layer2_outputs(9001)) xor (layer2_outputs(4135));
    outputs(7) <= not(layer2_outputs(8034));
    outputs(8) <= layer2_outputs(8597);
    outputs(9) <= layer2_outputs(630);
    outputs(10) <= not(layer2_outputs(2799));
    outputs(11) <= not(layer2_outputs(3492));
    outputs(12) <= layer2_outputs(100);
    outputs(13) <= not(layer2_outputs(8917));
    outputs(14) <= not((layer2_outputs(3788)) xor (layer2_outputs(4570)));
    outputs(15) <= not((layer2_outputs(1991)) xor (layer2_outputs(7214)));
    outputs(16) <= not(layer2_outputs(545));
    outputs(17) <= not(layer2_outputs(330));
    outputs(18) <= layer2_outputs(1651);
    outputs(19) <= layer2_outputs(9983);
    outputs(20) <= not(layer2_outputs(8712));
    outputs(21) <= layer2_outputs(1404);
    outputs(22) <= (layer2_outputs(1434)) and (layer2_outputs(2126));
    outputs(23) <= layer2_outputs(2723);
    outputs(24) <= not((layer2_outputs(9957)) or (layer2_outputs(7964)));
    outputs(25) <= not(layer2_outputs(3181));
    outputs(26) <= (layer2_outputs(1138)) or (layer2_outputs(8457));
    outputs(27) <= (layer2_outputs(7321)) and not (layer2_outputs(7669));
    outputs(28) <= not(layer2_outputs(8883));
    outputs(29) <= not((layer2_outputs(1363)) xor (layer2_outputs(5138)));
    outputs(30) <= (layer2_outputs(10017)) and (layer2_outputs(1364));
    outputs(31) <= not(layer2_outputs(334));
    outputs(32) <= layer2_outputs(453);
    outputs(33) <= not((layer2_outputs(3366)) and (layer2_outputs(9823)));
    outputs(34) <= layer2_outputs(8148);
    outputs(35) <= not((layer2_outputs(10076)) xor (layer2_outputs(10013)));
    outputs(36) <= not(layer2_outputs(6260)) or (layer2_outputs(9127));
    outputs(37) <= not(layer2_outputs(9348));
    outputs(38) <= not(layer2_outputs(8962));
    outputs(39) <= layer2_outputs(6775);
    outputs(40) <= layer2_outputs(1441);
    outputs(41) <= not(layer2_outputs(3595));
    outputs(42) <= (layer2_outputs(1252)) and not (layer2_outputs(7567));
    outputs(43) <= not(layer2_outputs(9258)) or (layer2_outputs(6188));
    outputs(44) <= layer2_outputs(8078);
    outputs(45) <= (layer2_outputs(3111)) xor (layer2_outputs(8272));
    outputs(46) <= not(layer2_outputs(4608));
    outputs(47) <= layer2_outputs(1603);
    outputs(48) <= not((layer2_outputs(4913)) xor (layer2_outputs(3868)));
    outputs(49) <= not((layer2_outputs(2479)) xor (layer2_outputs(9767)));
    outputs(50) <= not(layer2_outputs(6077));
    outputs(51) <= not(layer2_outputs(3264));
    outputs(52) <= not(layer2_outputs(6141));
    outputs(53) <= not(layer2_outputs(1472));
    outputs(54) <= (layer2_outputs(7120)) and not (layer2_outputs(2432));
    outputs(55) <= (layer2_outputs(336)) and not (layer2_outputs(8525));
    outputs(56) <= layer2_outputs(8846);
    outputs(57) <= layer2_outputs(1467);
    outputs(58) <= (layer2_outputs(5127)) or (layer2_outputs(5986));
    outputs(59) <= layer2_outputs(6239);
    outputs(60) <= layer2_outputs(4675);
    outputs(61) <= not((layer2_outputs(5436)) xor (layer2_outputs(8129)));
    outputs(62) <= (layer2_outputs(9226)) or (layer2_outputs(1654));
    outputs(63) <= not(layer2_outputs(2563)) or (layer2_outputs(5517));
    outputs(64) <= not((layer2_outputs(6399)) xor (layer2_outputs(4527)));
    outputs(65) <= layer2_outputs(3549);
    outputs(66) <= layer2_outputs(6436);
    outputs(67) <= not((layer2_outputs(6428)) xor (layer2_outputs(4245)));
    outputs(68) <= not(layer2_outputs(4959));
    outputs(69) <= not(layer2_outputs(10227)) or (layer2_outputs(9673));
    outputs(70) <= (layer2_outputs(5458)) and not (layer2_outputs(2120));
    outputs(71) <= (layer2_outputs(5873)) xor (layer2_outputs(2980));
    outputs(72) <= layer2_outputs(4019);
    outputs(73) <= not((layer2_outputs(3340)) xor (layer2_outputs(7936)));
    outputs(74) <= (layer2_outputs(5612)) xor (layer2_outputs(143));
    outputs(75) <= not(layer2_outputs(4855));
    outputs(76) <= layer2_outputs(7692);
    outputs(77) <= not(layer2_outputs(4234));
    outputs(78) <= (layer2_outputs(10200)) xor (layer2_outputs(9471));
    outputs(79) <= layer2_outputs(6179);
    outputs(80) <= not((layer2_outputs(5438)) or (layer2_outputs(5671)));
    outputs(81) <= not(layer2_outputs(553)) or (layer2_outputs(6331));
    outputs(82) <= not(layer2_outputs(6716));
    outputs(83) <= (layer2_outputs(5722)) or (layer2_outputs(3048));
    outputs(84) <= not(layer2_outputs(1029));
    outputs(85) <= (layer2_outputs(5955)) and not (layer2_outputs(5901));
    outputs(86) <= not(layer2_outputs(5768));
    outputs(87) <= not(layer2_outputs(4800));
    outputs(88) <= (layer2_outputs(8762)) xor (layer2_outputs(2013));
    outputs(89) <= not(layer2_outputs(1686)) or (layer2_outputs(321));
    outputs(90) <= not((layer2_outputs(5586)) or (layer2_outputs(3238)));
    outputs(91) <= layer2_outputs(7633);
    outputs(92) <= (layer2_outputs(3980)) xor (layer2_outputs(5636));
    outputs(93) <= not((layer2_outputs(9749)) xor (layer2_outputs(6161)));
    outputs(94) <= layer2_outputs(7828);
    outputs(95) <= layer2_outputs(943);
    outputs(96) <= layer2_outputs(2064);
    outputs(97) <= not(layer2_outputs(2309));
    outputs(98) <= not((layer2_outputs(491)) xor (layer2_outputs(211)));
    outputs(99) <= layer2_outputs(3894);
    outputs(100) <= (layer2_outputs(5612)) or (layer2_outputs(7684));
    outputs(101) <= (layer2_outputs(2452)) and (layer2_outputs(5490));
    outputs(102) <= layer2_outputs(904);
    outputs(103) <= not(layer2_outputs(10));
    outputs(104) <= not((layer2_outputs(7007)) or (layer2_outputs(4015)));
    outputs(105) <= not((layer2_outputs(2085)) xor (layer2_outputs(3877)));
    outputs(106) <= layer2_outputs(10225);
    outputs(107) <= layer2_outputs(2942);
    outputs(108) <= (layer2_outputs(2481)) and (layer2_outputs(1334));
    outputs(109) <= not(layer2_outputs(6600));
    outputs(110) <= layer2_outputs(8957);
    outputs(111) <= not((layer2_outputs(4146)) xor (layer2_outputs(2798)));
    outputs(112) <= not(layer2_outputs(4139));
    outputs(113) <= not(layer2_outputs(1874));
    outputs(114) <= (layer2_outputs(5889)) xor (layer2_outputs(519));
    outputs(115) <= not(layer2_outputs(6909)) or (layer2_outputs(10072));
    outputs(116) <= not(layer2_outputs(8747)) or (layer2_outputs(4216));
    outputs(117) <= (layer2_outputs(2004)) xor (layer2_outputs(7433));
    outputs(118) <= (layer2_outputs(211)) and (layer2_outputs(4481));
    outputs(119) <= (layer2_outputs(9962)) and not (layer2_outputs(9442));
    outputs(120) <= layer2_outputs(4721);
    outputs(121) <= not(layer2_outputs(7294));
    outputs(122) <= layer2_outputs(5625);
    outputs(123) <= layer2_outputs(1280);
    outputs(124) <= layer2_outputs(1314);
    outputs(125) <= not(layer2_outputs(9988));
    outputs(126) <= (layer2_outputs(9670)) and not (layer2_outputs(8817));
    outputs(127) <= (layer2_outputs(1752)) or (layer2_outputs(3945));
    outputs(128) <= not(layer2_outputs(6198));
    outputs(129) <= not(layer2_outputs(7485));
    outputs(130) <= not((layer2_outputs(1938)) or (layer2_outputs(67)));
    outputs(131) <= layer2_outputs(18);
    outputs(132) <= not((layer2_outputs(3077)) or (layer2_outputs(7510)));
    outputs(133) <= not((layer2_outputs(6662)) xor (layer2_outputs(10236)));
    outputs(134) <= not((layer2_outputs(4801)) xor (layer2_outputs(2028)));
    outputs(135) <= not(layer2_outputs(5371));
    outputs(136) <= not(layer2_outputs(5400));
    outputs(137) <= layer2_outputs(6960);
    outputs(138) <= layer2_outputs(10049);
    outputs(139) <= not(layer2_outputs(8476));
    outputs(140) <= (layer2_outputs(423)) and not (layer2_outputs(7119));
    outputs(141) <= not(layer2_outputs(89));
    outputs(142) <= (layer2_outputs(2129)) xor (layer2_outputs(2691));
    outputs(143) <= not(layer2_outputs(9514));
    outputs(144) <= (layer2_outputs(1091)) and (layer2_outputs(7993));
    outputs(145) <= not(layer2_outputs(2196));
    outputs(146) <= not(layer2_outputs(5039));
    outputs(147) <= (layer2_outputs(6591)) xor (layer2_outputs(5984));
    outputs(148) <= layer2_outputs(4593);
    outputs(149) <= layer2_outputs(1272);
    outputs(150) <= layer2_outputs(3355);
    outputs(151) <= (layer2_outputs(186)) xor (layer2_outputs(6545));
    outputs(152) <= not((layer2_outputs(1128)) xor (layer2_outputs(3984)));
    outputs(153) <= not(layer2_outputs(2409));
    outputs(154) <= layer2_outputs(9454);
    outputs(155) <= not((layer2_outputs(3626)) xor (layer2_outputs(2774)));
    outputs(156) <= (layer2_outputs(6731)) xor (layer2_outputs(6126));
    outputs(157) <= (layer2_outputs(2283)) and (layer2_outputs(6185));
    outputs(158) <= not((layer2_outputs(6356)) xor (layer2_outputs(6197)));
    outputs(159) <= not(layer2_outputs(3370));
    outputs(160) <= not(layer2_outputs(9622));
    outputs(161) <= not(layer2_outputs(1697));
    outputs(162) <= not(layer2_outputs(5003));
    outputs(163) <= (layer2_outputs(9406)) xor (layer2_outputs(10103));
    outputs(164) <= not(layer2_outputs(2276));
    outputs(165) <= (layer2_outputs(9343)) and not (layer2_outputs(7880));
    outputs(166) <= (layer2_outputs(8619)) and not (layer2_outputs(8247));
    outputs(167) <= (layer2_outputs(1161)) and (layer2_outputs(9502));
    outputs(168) <= (layer2_outputs(8377)) and not (layer2_outputs(2150));
    outputs(169) <= layer2_outputs(1993);
    outputs(170) <= layer2_outputs(5);
    outputs(171) <= not(layer2_outputs(9258));
    outputs(172) <= layer2_outputs(5894);
    outputs(173) <= (layer2_outputs(1078)) or (layer2_outputs(10022));
    outputs(174) <= not(layer2_outputs(9189));
    outputs(175) <= not(layer2_outputs(8381));
    outputs(176) <= not(layer2_outputs(6447));
    outputs(177) <= layer2_outputs(2056);
    outputs(178) <= layer2_outputs(6461);
    outputs(179) <= (layer2_outputs(5268)) or (layer2_outputs(9058));
    outputs(180) <= layer2_outputs(7335);
    outputs(181) <= not(layer2_outputs(9643));
    outputs(182) <= not((layer2_outputs(9165)) xor (layer2_outputs(2762)));
    outputs(183) <= layer2_outputs(4386);
    outputs(184) <= (layer2_outputs(7200)) and (layer2_outputs(332));
    outputs(185) <= (layer2_outputs(5685)) and not (layer2_outputs(4960));
    outputs(186) <= not(layer2_outputs(564));
    outputs(187) <= not(layer2_outputs(4053));
    outputs(188) <= not((layer2_outputs(1709)) xor (layer2_outputs(9833)));
    outputs(189) <= layer2_outputs(1481);
    outputs(190) <= (layer2_outputs(3605)) and not (layer2_outputs(5344));
    outputs(191) <= not(layer2_outputs(5640));
    outputs(192) <= layer2_outputs(5146);
    outputs(193) <= layer2_outputs(7751);
    outputs(194) <= layer2_outputs(7272);
    outputs(195) <= not((layer2_outputs(5569)) or (layer2_outputs(1356)));
    outputs(196) <= (layer2_outputs(3119)) and not (layer2_outputs(2432));
    outputs(197) <= not(layer2_outputs(7062));
    outputs(198) <= layer2_outputs(3630);
    outputs(199) <= (layer2_outputs(150)) and not (layer2_outputs(5702));
    outputs(200) <= layer2_outputs(4490);
    outputs(201) <= layer2_outputs(100);
    outputs(202) <= layer2_outputs(6165);
    outputs(203) <= layer2_outputs(2530);
    outputs(204) <= layer2_outputs(6062);
    outputs(205) <= not(layer2_outputs(8114));
    outputs(206) <= not((layer2_outputs(1869)) xor (layer2_outputs(1587)));
    outputs(207) <= layer2_outputs(604);
    outputs(208) <= layer2_outputs(8834);
    outputs(209) <= layer2_outputs(3332);
    outputs(210) <= (layer2_outputs(3133)) xor (layer2_outputs(3149));
    outputs(211) <= (layer2_outputs(7743)) and not (layer2_outputs(5134));
    outputs(212) <= not((layer2_outputs(9270)) xor (layer2_outputs(2649)));
    outputs(213) <= layer2_outputs(8233);
    outputs(214) <= not(layer2_outputs(6947));
    outputs(215) <= not(layer2_outputs(441));
    outputs(216) <= not(layer2_outputs(4152));
    outputs(217) <= layer2_outputs(6702);
    outputs(218) <= (layer2_outputs(2082)) xor (layer2_outputs(496));
    outputs(219) <= not((layer2_outputs(7091)) xor (layer2_outputs(547)));
    outputs(220) <= not((layer2_outputs(5473)) or (layer2_outputs(514)));
    outputs(221) <= not(layer2_outputs(611)) or (layer2_outputs(4286));
    outputs(222) <= not((layer2_outputs(4661)) and (layer2_outputs(3817)));
    outputs(223) <= (layer2_outputs(3246)) and (layer2_outputs(1649));
    outputs(224) <= layer2_outputs(7744);
    outputs(225) <= (layer2_outputs(7260)) xor (layer2_outputs(4117));
    outputs(226) <= not(layer2_outputs(3834)) or (layer2_outputs(7262));
    outputs(227) <= not((layer2_outputs(9877)) xor (layer2_outputs(8029)));
    outputs(228) <= not(layer2_outputs(6057));
    outputs(229) <= (layer2_outputs(5590)) or (layer2_outputs(1024));
    outputs(230) <= (layer2_outputs(2606)) xor (layer2_outputs(8759));
    outputs(231) <= not(layer2_outputs(3190));
    outputs(232) <= not(layer2_outputs(2795));
    outputs(233) <= (layer2_outputs(8487)) xor (layer2_outputs(2759));
    outputs(234) <= layer2_outputs(2428);
    outputs(235) <= layer2_outputs(3221);
    outputs(236) <= (layer2_outputs(9188)) and not (layer2_outputs(7990));
    outputs(237) <= (layer2_outputs(38)) and not (layer2_outputs(9808));
    outputs(238) <= layer2_outputs(2324);
    outputs(239) <= layer2_outputs(8665);
    outputs(240) <= layer2_outputs(787);
    outputs(241) <= (layer2_outputs(366)) xor (layer2_outputs(6362));
    outputs(242) <= not((layer2_outputs(9156)) or (layer2_outputs(2768)));
    outputs(243) <= not(layer2_outputs(340));
    outputs(244) <= not(layer2_outputs(1388));
    outputs(245) <= not(layer2_outputs(9665));
    outputs(246) <= not(layer2_outputs(852));
    outputs(247) <= (layer2_outputs(7752)) and not (layer2_outputs(6360));
    outputs(248) <= layer2_outputs(1689);
    outputs(249) <= layer2_outputs(6615);
    outputs(250) <= not(layer2_outputs(9509));
    outputs(251) <= not(layer2_outputs(507));
    outputs(252) <= (layer2_outputs(2062)) and not (layer2_outputs(5324));
    outputs(253) <= layer2_outputs(9828);
    outputs(254) <= not((layer2_outputs(3633)) or (layer2_outputs(5036)));
    outputs(255) <= layer2_outputs(1811);
    outputs(256) <= (layer2_outputs(7287)) and not (layer2_outputs(9234));
    outputs(257) <= not((layer2_outputs(3778)) xor (layer2_outputs(1342)));
    outputs(258) <= not(layer2_outputs(7578));
    outputs(259) <= not((layer2_outputs(8111)) or (layer2_outputs(3573)));
    outputs(260) <= (layer2_outputs(7786)) and (layer2_outputs(1039));
    outputs(261) <= (layer2_outputs(1271)) xor (layer2_outputs(9676));
    outputs(262) <= layer2_outputs(8442);
    outputs(263) <= not(layer2_outputs(2841)) or (layer2_outputs(108));
    outputs(264) <= not(layer2_outputs(4987)) or (layer2_outputs(7045));
    outputs(265) <= layer2_outputs(1014);
    outputs(266) <= (layer2_outputs(1306)) and not (layer2_outputs(1462));
    outputs(267) <= not(layer2_outputs(7625));
    outputs(268) <= not((layer2_outputs(9794)) or (layer2_outputs(1624)));
    outputs(269) <= not((layer2_outputs(7172)) and (layer2_outputs(8870)));
    outputs(270) <= not(layer2_outputs(3197)) or (layer2_outputs(8241));
    outputs(271) <= not((layer2_outputs(886)) xor (layer2_outputs(2425)));
    outputs(272) <= layer2_outputs(5531);
    outputs(273) <= not(layer2_outputs(8098));
    outputs(274) <= not((layer2_outputs(4957)) xor (layer2_outputs(3855)));
    outputs(275) <= not(layer2_outputs(51));
    outputs(276) <= (layer2_outputs(6743)) and not (layer2_outputs(653));
    outputs(277) <= not(layer2_outputs(5377));
    outputs(278) <= (layer2_outputs(1926)) xor (layer2_outputs(8774));
    outputs(279) <= layer2_outputs(1671);
    outputs(280) <= not(layer2_outputs(3209)) or (layer2_outputs(8236));
    outputs(281) <= (layer2_outputs(9530)) and not (layer2_outputs(5887));
    outputs(282) <= not(layer2_outputs(6554)) or (layer2_outputs(7965));
    outputs(283) <= not(layer2_outputs(4013));
    outputs(284) <= not(layer2_outputs(8543));
    outputs(285) <= not(layer2_outputs(5449)) or (layer2_outputs(9559));
    outputs(286) <= layer2_outputs(2724);
    outputs(287) <= not(layer2_outputs(7386));
    outputs(288) <= layer2_outputs(4176);
    outputs(289) <= layer2_outputs(9510);
    outputs(290) <= layer2_outputs(2542);
    outputs(291) <= not(layer2_outputs(6233));
    outputs(292) <= not((layer2_outputs(6155)) and (layer2_outputs(5264)));
    outputs(293) <= layer2_outputs(9082);
    outputs(294) <= not(layer2_outputs(5707));
    outputs(295) <= (layer2_outputs(244)) or (layer2_outputs(7270));
    outputs(296) <= not(layer2_outputs(596));
    outputs(297) <= not(layer2_outputs(4620));
    outputs(298) <= not(layer2_outputs(7622));
    outputs(299) <= not(layer2_outputs(8892)) or (layer2_outputs(741));
    outputs(300) <= not(layer2_outputs(5008));
    outputs(301) <= layer2_outputs(10222);
    outputs(302) <= not((layer2_outputs(371)) and (layer2_outputs(8410)));
    outputs(303) <= not(layer2_outputs(5061));
    outputs(304) <= layer2_outputs(2901);
    outputs(305) <= layer2_outputs(6551);
    outputs(306) <= not((layer2_outputs(7142)) or (layer2_outputs(1230)));
    outputs(307) <= not((layer2_outputs(6375)) xor (layer2_outputs(9231)));
    outputs(308) <= layer2_outputs(3270);
    outputs(309) <= layer2_outputs(2512);
    outputs(310) <= not(layer2_outputs(3783));
    outputs(311) <= layer2_outputs(4204);
    outputs(312) <= not(layer2_outputs(7244));
    outputs(313) <= not(layer2_outputs(4793));
    outputs(314) <= layer2_outputs(3171);
    outputs(315) <= layer2_outputs(3620);
    outputs(316) <= layer2_outputs(6992);
    outputs(317) <= not((layer2_outputs(8312)) or (layer2_outputs(3673)));
    outputs(318) <= layer2_outputs(5995);
    outputs(319) <= layer2_outputs(2173);
    outputs(320) <= layer2_outputs(1319);
    outputs(321) <= layer2_outputs(2491);
    outputs(322) <= layer2_outputs(2891);
    outputs(323) <= not((layer2_outputs(6402)) xor (layer2_outputs(2564)));
    outputs(324) <= layer2_outputs(642);
    outputs(325) <= (layer2_outputs(4689)) xor (layer2_outputs(4816));
    outputs(326) <= not(layer2_outputs(3923));
    outputs(327) <= not(layer2_outputs(3636));
    outputs(328) <= layer2_outputs(8308);
    outputs(329) <= layer2_outputs(8182);
    outputs(330) <= layer2_outputs(6881);
    outputs(331) <= layer2_outputs(1481);
    outputs(332) <= (layer2_outputs(6124)) or (layer2_outputs(8355));
    outputs(333) <= not(layer2_outputs(3981));
    outputs(334) <= not(layer2_outputs(5335));
    outputs(335) <= not(layer2_outputs(1249));
    outputs(336) <= layer2_outputs(7399);
    outputs(337) <= layer2_outputs(7263);
    outputs(338) <= (layer2_outputs(7044)) and not (layer2_outputs(5219));
    outputs(339) <= layer2_outputs(910);
    outputs(340) <= layer2_outputs(5112);
    outputs(341) <= (layer2_outputs(6081)) xor (layer2_outputs(333));
    outputs(342) <= not((layer2_outputs(2665)) xor (layer2_outputs(2482)));
    outputs(343) <= not(layer2_outputs(3418));
    outputs(344) <= layer2_outputs(1853);
    outputs(345) <= not(layer2_outputs(5372));
    outputs(346) <= layer2_outputs(8545);
    outputs(347) <= not(layer2_outputs(8794));
    outputs(348) <= layer2_outputs(3836);
    outputs(349) <= (layer2_outputs(3271)) and (layer2_outputs(4555));
    outputs(350) <= not((layer2_outputs(1848)) xor (layer2_outputs(3465)));
    outputs(351) <= layer2_outputs(9534);
    outputs(352) <= layer2_outputs(1925);
    outputs(353) <= not(layer2_outputs(8306));
    outputs(354) <= layer2_outputs(372);
    outputs(355) <= (layer2_outputs(2630)) xor (layer2_outputs(6345));
    outputs(356) <= layer2_outputs(85);
    outputs(357) <= layer2_outputs(7712);
    outputs(358) <= (layer2_outputs(768)) xor (layer2_outputs(4216));
    outputs(359) <= layer2_outputs(7916);
    outputs(360) <= not(layer2_outputs(7145)) or (layer2_outputs(4943));
    outputs(361) <= layer2_outputs(5498);
    outputs(362) <= not((layer2_outputs(2356)) xor (layer2_outputs(8235)));
    outputs(363) <= (layer2_outputs(5630)) and (layer2_outputs(6347));
    outputs(364) <= layer2_outputs(5293);
    outputs(365) <= layer2_outputs(65);
    outputs(366) <= (layer2_outputs(3277)) and not (layer2_outputs(555));
    outputs(367) <= (layer2_outputs(4867)) or (layer2_outputs(4425));
    outputs(368) <= not(layer2_outputs(9293));
    outputs(369) <= (layer2_outputs(2066)) xor (layer2_outputs(3700));
    outputs(370) <= layer2_outputs(4879);
    outputs(371) <= layer2_outputs(3329);
    outputs(372) <= not(layer2_outputs(2662));
    outputs(373) <= layer2_outputs(2610);
    outputs(374) <= layer2_outputs(1638);
    outputs(375) <= layer2_outputs(6291);
    outputs(376) <= layer2_outputs(4632);
    outputs(377) <= not(layer2_outputs(8486));
    outputs(378) <= (layer2_outputs(8984)) xor (layer2_outputs(212));
    outputs(379) <= not(layer2_outputs(6039));
    outputs(380) <= layer2_outputs(4796);
    outputs(381) <= not(layer2_outputs(7593));
    outputs(382) <= (layer2_outputs(4918)) or (layer2_outputs(2506));
    outputs(383) <= not(layer2_outputs(10216));
    outputs(384) <= not(layer2_outputs(2496));
    outputs(385) <= (layer2_outputs(10090)) xor (layer2_outputs(1267));
    outputs(386) <= not(layer2_outputs(6205));
    outputs(387) <= not(layer2_outputs(7708));
    outputs(388) <= layer2_outputs(1967);
    outputs(389) <= not(layer2_outputs(3815));
    outputs(390) <= layer2_outputs(4020);
    outputs(391) <= (layer2_outputs(8446)) and not (layer2_outputs(7589));
    outputs(392) <= not(layer2_outputs(535));
    outputs(393) <= not((layer2_outputs(8803)) xor (layer2_outputs(3748)));
    outputs(394) <= layer2_outputs(639);
    outputs(395) <= layer2_outputs(4442);
    outputs(396) <= (layer2_outputs(10155)) and (layer2_outputs(7775));
    outputs(397) <= not((layer2_outputs(8955)) or (layer2_outputs(6953)));
    outputs(398) <= (layer2_outputs(4580)) and (layer2_outputs(3763));
    outputs(399) <= (layer2_outputs(4257)) and not (layer2_outputs(5906));
    outputs(400) <= layer2_outputs(3609);
    outputs(401) <= layer2_outputs(7734);
    outputs(402) <= layer2_outputs(9109);
    outputs(403) <= not(layer2_outputs(2247));
    outputs(404) <= layer2_outputs(5118);
    outputs(405) <= layer2_outputs(1143);
    outputs(406) <= layer2_outputs(6522);
    outputs(407) <= layer2_outputs(999);
    outputs(408) <= layer2_outputs(7381);
    outputs(409) <= not(layer2_outputs(4269));
    outputs(410) <= layer2_outputs(8483);
    outputs(411) <= not((layer2_outputs(9420)) xor (layer2_outputs(8277)));
    outputs(412) <= layer2_outputs(8196);
    outputs(413) <= not((layer2_outputs(2726)) and (layer2_outputs(7172)));
    outputs(414) <= not(layer2_outputs(3557));
    outputs(415) <= not((layer2_outputs(7976)) xor (layer2_outputs(3109)));
    outputs(416) <= (layer2_outputs(9286)) xor (layer2_outputs(9486));
    outputs(417) <= not(layer2_outputs(8114)) or (layer2_outputs(1486));
    outputs(418) <= not((layer2_outputs(9289)) xor (layer2_outputs(7031)));
    outputs(419) <= not(layer2_outputs(5257));
    outputs(420) <= layer2_outputs(483);
    outputs(421) <= not((layer2_outputs(255)) xor (layer2_outputs(1245)));
    outputs(422) <= (layer2_outputs(6824)) xor (layer2_outputs(1025));
    outputs(423) <= not(layer2_outputs(797));
    outputs(424) <= not(layer2_outputs(5488)) or (layer2_outputs(4411));
    outputs(425) <= layer2_outputs(1988);
    outputs(426) <= layer2_outputs(5091);
    outputs(427) <= layer2_outputs(1458);
    outputs(428) <= not(layer2_outputs(5818)) or (layer2_outputs(7313));
    outputs(429) <= layer2_outputs(489);
    outputs(430) <= not(layer2_outputs(949));
    outputs(431) <= not((layer2_outputs(2934)) and (layer2_outputs(8731)));
    outputs(432) <= not(layer2_outputs(9151));
    outputs(433) <= layer2_outputs(5441);
    outputs(434) <= (layer2_outputs(993)) xor (layer2_outputs(3631));
    outputs(435) <= not((layer2_outputs(8713)) xor (layer2_outputs(7428)));
    outputs(436) <= not(layer2_outputs(5953)) or (layer2_outputs(8707));
    outputs(437) <= not(layer2_outputs(685));
    outputs(438) <= not(layer2_outputs(7286)) or (layer2_outputs(9673));
    outputs(439) <= not((layer2_outputs(656)) xor (layer2_outputs(7443)));
    outputs(440) <= (layer2_outputs(4129)) xor (layer2_outputs(4552));
    outputs(441) <= layer2_outputs(2637);
    outputs(442) <= not(layer2_outputs(9218));
    outputs(443) <= not(layer2_outputs(4747));
    outputs(444) <= layer2_outputs(630);
    outputs(445) <= not(layer2_outputs(3681));
    outputs(446) <= (layer2_outputs(2221)) and not (layer2_outputs(7726));
    outputs(447) <= not(layer2_outputs(2742));
    outputs(448) <= layer2_outputs(4002);
    outputs(449) <= not((layer2_outputs(7652)) xor (layer2_outputs(2508)));
    outputs(450) <= (layer2_outputs(4885)) and not (layer2_outputs(3946));
    outputs(451) <= layer2_outputs(6815);
    outputs(452) <= not(layer2_outputs(661));
    outputs(453) <= not(layer2_outputs(9055));
    outputs(454) <= not(layer2_outputs(1211));
    outputs(455) <= not(layer2_outputs(6949));
    outputs(456) <= not((layer2_outputs(8324)) xor (layer2_outputs(4138)));
    outputs(457) <= not(layer2_outputs(4344));
    outputs(458) <= not(layer2_outputs(1827));
    outputs(459) <= not((layer2_outputs(6950)) xor (layer2_outputs(7148)));
    outputs(460) <= not((layer2_outputs(10164)) xor (layer2_outputs(9915)));
    outputs(461) <= not((layer2_outputs(407)) xor (layer2_outputs(2504)));
    outputs(462) <= not(layer2_outputs(9080));
    outputs(463) <= layer2_outputs(7012);
    outputs(464) <= not((layer2_outputs(3434)) and (layer2_outputs(9363)));
    outputs(465) <= (layer2_outputs(7526)) xor (layer2_outputs(4285));
    outputs(466) <= (layer2_outputs(4754)) and not (layer2_outputs(4479));
    outputs(467) <= not((layer2_outputs(10036)) or (layer2_outputs(4601)));
    outputs(468) <= layer2_outputs(7317);
    outputs(469) <= not(layer2_outputs(3406));
    outputs(470) <= not(layer2_outputs(8455));
    outputs(471) <= not(layer2_outputs(2195));
    outputs(472) <= not((layer2_outputs(3775)) xor (layer2_outputs(307)));
    outputs(473) <= layer2_outputs(7986);
    outputs(474) <= not(layer2_outputs(7973));
    outputs(475) <= not(layer2_outputs(3244));
    outputs(476) <= (layer2_outputs(8230)) and not (layer2_outputs(5952));
    outputs(477) <= not(layer2_outputs(4209));
    outputs(478) <= layer2_outputs(9317);
    outputs(479) <= layer2_outputs(2011);
    outputs(480) <= not(layer2_outputs(4051));
    outputs(481) <= layer2_outputs(2352);
    outputs(482) <= layer2_outputs(6423);
    outputs(483) <= (layer2_outputs(5823)) and not (layer2_outputs(9985));
    outputs(484) <= not(layer2_outputs(7803)) or (layer2_outputs(3004));
    outputs(485) <= not(layer2_outputs(2147));
    outputs(486) <= (layer2_outputs(882)) and not (layer2_outputs(2547));
    outputs(487) <= not(layer2_outputs(4041));
    outputs(488) <= (layer2_outputs(3581)) or (layer2_outputs(1259));
    outputs(489) <= layer2_outputs(251);
    outputs(490) <= layer2_outputs(9777);
    outputs(491) <= (layer2_outputs(1117)) and not (layer2_outputs(7943));
    outputs(492) <= not((layer2_outputs(2785)) xor (layer2_outputs(4450)));
    outputs(493) <= (layer2_outputs(9685)) and not (layer2_outputs(4008));
    outputs(494) <= layer2_outputs(7674);
    outputs(495) <= not((layer2_outputs(8433)) xor (layer2_outputs(3408)));
    outputs(496) <= not(layer2_outputs(2771));
    outputs(497) <= not(layer2_outputs(12));
    outputs(498) <= (layer2_outputs(8931)) xor (layer2_outputs(68));
    outputs(499) <= not((layer2_outputs(6978)) xor (layer2_outputs(6439)));
    outputs(500) <= layer2_outputs(149);
    outputs(501) <= not((layer2_outputs(6576)) xor (layer2_outputs(5747)));
    outputs(502) <= (layer2_outputs(55)) and not (layer2_outputs(9711));
    outputs(503) <= layer2_outputs(608);
    outputs(504) <= (layer2_outputs(2800)) and not (layer2_outputs(2347));
    outputs(505) <= layer2_outputs(3410);
    outputs(506) <= layer2_outputs(6247);
    outputs(507) <= (layer2_outputs(9096)) and not (layer2_outputs(1681));
    outputs(508) <= layer2_outputs(2578);
    outputs(509) <= not(layer2_outputs(3591));
    outputs(510) <= layer2_outputs(2045);
    outputs(511) <= layer2_outputs(7497);
    outputs(512) <= (layer2_outputs(2943)) xor (layer2_outputs(6973));
    outputs(513) <= not(layer2_outputs(5399));
    outputs(514) <= layer2_outputs(4487);
    outputs(515) <= not((layer2_outputs(3904)) xor (layer2_outputs(6635)));
    outputs(516) <= (layer2_outputs(7047)) and not (layer2_outputs(2300));
    outputs(517) <= layer2_outputs(733);
    outputs(518) <= layer2_outputs(2894);
    outputs(519) <= not(layer2_outputs(8430));
    outputs(520) <= layer2_outputs(7125);
    outputs(521) <= layer2_outputs(3995);
    outputs(522) <= not((layer2_outputs(9615)) and (layer2_outputs(9168)));
    outputs(523) <= not(layer2_outputs(5998));
    outputs(524) <= not((layer2_outputs(599)) xor (layer2_outputs(2488)));
    outputs(525) <= (layer2_outputs(2887)) and not (layer2_outputs(1665));
    outputs(526) <= not(layer2_outputs(9799));
    outputs(527) <= not(layer2_outputs(2255));
    outputs(528) <= layer2_outputs(3786);
    outputs(529) <= layer2_outputs(680);
    outputs(530) <= not(layer2_outputs(626));
    outputs(531) <= not((layer2_outputs(6324)) or (layer2_outputs(5252)));
    outputs(532) <= (layer2_outputs(6907)) and (layer2_outputs(5237));
    outputs(533) <= layer2_outputs(2543);
    outputs(534) <= (layer2_outputs(6819)) xor (layer2_outputs(6425));
    outputs(535) <= not(layer2_outputs(3458)) or (layer2_outputs(5247));
    outputs(536) <= not(layer2_outputs(7388));
    outputs(537) <= (layer2_outputs(1419)) xor (layer2_outputs(4915));
    outputs(538) <= not(layer2_outputs(9390));
    outputs(539) <= not(layer2_outputs(6984));
    outputs(540) <= layer2_outputs(4714);
    outputs(541) <= not(layer2_outputs(2613));
    outputs(542) <= not(layer2_outputs(6498)) or (layer2_outputs(9633));
    outputs(543) <= layer2_outputs(8601);
    outputs(544) <= layer2_outputs(2610);
    outputs(545) <= not(layer2_outputs(7689));
    outputs(546) <= not(layer2_outputs(4963));
    outputs(547) <= layer2_outputs(6812);
    outputs(548) <= (layer2_outputs(913)) xor (layer2_outputs(1947));
    outputs(549) <= not(layer2_outputs(6311));
    outputs(550) <= (layer2_outputs(7781)) xor (layer2_outputs(4341));
    outputs(551) <= not((layer2_outputs(58)) and (layer2_outputs(815)));
    outputs(552) <= (layer2_outputs(3230)) xor (layer2_outputs(9391));
    outputs(553) <= layer2_outputs(7283);
    outputs(554) <= (layer2_outputs(1719)) and not (layer2_outputs(3005));
    outputs(555) <= not((layer2_outputs(8687)) and (layer2_outputs(9574)));
    outputs(556) <= (layer2_outputs(9328)) xor (layer2_outputs(4606));
    outputs(557) <= not((layer2_outputs(8543)) or (layer2_outputs(6774)));
    outputs(558) <= layer2_outputs(9056);
    outputs(559) <= not(layer2_outputs(5710));
    outputs(560) <= (layer2_outputs(5062)) and (layer2_outputs(3262));
    outputs(561) <= not((layer2_outputs(9573)) xor (layer2_outputs(7032)));
    outputs(562) <= not(layer2_outputs(6685));
    outputs(563) <= (layer2_outputs(625)) and not (layer2_outputs(1125));
    outputs(564) <= not(layer2_outputs(7147)) or (layer2_outputs(5938));
    outputs(565) <= not(layer2_outputs(10218));
    outputs(566) <= layer2_outputs(8649);
    outputs(567) <= not(layer2_outputs(9040));
    outputs(568) <= layer2_outputs(5173);
    outputs(569) <= not((layer2_outputs(1741)) or (layer2_outputs(4670)));
    outputs(570) <= not(layer2_outputs(2749));
    outputs(571) <= layer2_outputs(5185);
    outputs(572) <= not(layer2_outputs(2052));
    outputs(573) <= (layer2_outputs(9621)) and not (layer2_outputs(2574));
    outputs(574) <= (layer2_outputs(3405)) or (layer2_outputs(1012));
    outputs(575) <= layer2_outputs(1621);
    outputs(576) <= not(layer2_outputs(7258));
    outputs(577) <= not(layer2_outputs(7232));
    outputs(578) <= layer2_outputs(10049);
    outputs(579) <= not((layer2_outputs(2738)) or (layer2_outputs(2255)));
    outputs(580) <= not(layer2_outputs(1738));
    outputs(581) <= not((layer2_outputs(3746)) or (layer2_outputs(545)));
    outputs(582) <= layer2_outputs(6013);
    outputs(583) <= not((layer2_outputs(5975)) xor (layer2_outputs(2715)));
    outputs(584) <= layer2_outputs(9157);
    outputs(585) <= layer2_outputs(4164);
    outputs(586) <= not((layer2_outputs(7006)) xor (layer2_outputs(5227)));
    outputs(587) <= layer2_outputs(1604);
    outputs(588) <= (layer2_outputs(9141)) and not (layer2_outputs(5989));
    outputs(589) <= (layer2_outputs(674)) xor (layer2_outputs(2042));
    outputs(590) <= layer2_outputs(5802);
    outputs(591) <= layer2_outputs(9109);
    outputs(592) <= not((layer2_outputs(2273)) or (layer2_outputs(7087)));
    outputs(593) <= not(layer2_outputs(6925));
    outputs(594) <= (layer2_outputs(7619)) and (layer2_outputs(7897));
    outputs(595) <= not(layer2_outputs(3696));
    outputs(596) <= not((layer2_outputs(648)) or (layer2_outputs(4631)));
    outputs(597) <= not(layer2_outputs(4273));
    outputs(598) <= layer2_outputs(8342);
    outputs(599) <= (layer2_outputs(1399)) and not (layer2_outputs(988));
    outputs(600) <= layer2_outputs(9096);
    outputs(601) <= not((layer2_outputs(2685)) xor (layer2_outputs(627)));
    outputs(602) <= not(layer2_outputs(74));
    outputs(603) <= not(layer2_outputs(8512));
    outputs(604) <= (layer2_outputs(6285)) and (layer2_outputs(5368));
    outputs(605) <= not((layer2_outputs(10133)) or (layer2_outputs(795)));
    outputs(606) <= (layer2_outputs(7512)) xor (layer2_outputs(285));
    outputs(607) <= (layer2_outputs(5791)) xor (layer2_outputs(2436));
    outputs(608) <= not(layer2_outputs(341));
    outputs(609) <= layer2_outputs(779);
    outputs(610) <= layer2_outputs(702);
    outputs(611) <= not(layer2_outputs(1483));
    outputs(612) <= (layer2_outputs(4971)) and (layer2_outputs(2769));
    outputs(613) <= not(layer2_outputs(5269)) or (layer2_outputs(6825));
    outputs(614) <= (layer2_outputs(8338)) xor (layer2_outputs(7693));
    outputs(615) <= layer2_outputs(7736);
    outputs(616) <= layer2_outputs(4627);
    outputs(617) <= layer2_outputs(138);
    outputs(618) <= (layer2_outputs(7030)) and not (layer2_outputs(970));
    outputs(619) <= layer2_outputs(4176);
    outputs(620) <= not(layer2_outputs(6206)) or (layer2_outputs(6759));
    outputs(621) <= (layer2_outputs(5742)) and not (layer2_outputs(4403));
    outputs(622) <= layer2_outputs(9922);
    outputs(623) <= layer2_outputs(4312);
    outputs(624) <= (layer2_outputs(5655)) and not (layer2_outputs(461));
    outputs(625) <= (layer2_outputs(6438)) and not (layer2_outputs(4447));
    outputs(626) <= layer2_outputs(2839);
    outputs(627) <= not(layer2_outputs(1432));
    outputs(628) <= not(layer2_outputs(2393)) or (layer2_outputs(3713));
    outputs(629) <= layer2_outputs(6151);
    outputs(630) <= layer2_outputs(6330);
    outputs(631) <= (layer2_outputs(8422)) and (layer2_outputs(4572));
    outputs(632) <= not((layer2_outputs(6282)) xor (layer2_outputs(5453)));
    outputs(633) <= (layer2_outputs(5809)) and not (layer2_outputs(8403));
    outputs(634) <= not(layer2_outputs(6599)) or (layer2_outputs(549));
    outputs(635) <= not(layer2_outputs(1824));
    outputs(636) <= layer2_outputs(8675);
    outputs(637) <= layer2_outputs(8404);
    outputs(638) <= (layer2_outputs(1768)) xor (layer2_outputs(1199));
    outputs(639) <= layer2_outputs(8116);
    outputs(640) <= not(layer2_outputs(9988));
    outputs(641) <= (layer2_outputs(9004)) xor (layer2_outputs(3372));
    outputs(642) <= (layer2_outputs(2070)) and not (layer2_outputs(7783));
    outputs(643) <= not(layer2_outputs(5887));
    outputs(644) <= not(layer2_outputs(4980));
    outputs(645) <= not(layer2_outputs(6891)) or (layer2_outputs(9044));
    outputs(646) <= (layer2_outputs(10205)) and (layer2_outputs(1364));
    outputs(647) <= (layer2_outputs(6671)) and (layer2_outputs(2389));
    outputs(648) <= (layer2_outputs(3339)) and (layer2_outputs(9705));
    outputs(649) <= (layer2_outputs(6659)) and (layer2_outputs(7146));
    outputs(650) <= not(layer2_outputs(4089));
    outputs(651) <= not((layer2_outputs(2196)) and (layer2_outputs(9947)));
    outputs(652) <= (layer2_outputs(9330)) and not (layer2_outputs(6193));
    outputs(653) <= layer2_outputs(6148);
    outputs(654) <= (layer2_outputs(5929)) and (layer2_outputs(4408));
    outputs(655) <= layer2_outputs(4905);
    outputs(656) <= not((layer2_outputs(2046)) xor (layer2_outputs(5019)));
    outputs(657) <= not(layer2_outputs(8371));
    outputs(658) <= not(layer2_outputs(9280));
    outputs(659) <= layer2_outputs(3894);
    outputs(660) <= not((layer2_outputs(3636)) xor (layer2_outputs(191)));
    outputs(661) <= not(layer2_outputs(7315)) or (layer2_outputs(9884));
    outputs(662) <= not((layer2_outputs(9545)) or (layer2_outputs(9423)));
    outputs(663) <= layer2_outputs(5931);
    outputs(664) <= not(layer2_outputs(7198));
    outputs(665) <= layer2_outputs(633);
    outputs(666) <= not(layer2_outputs(2895));
    outputs(667) <= not(layer2_outputs(8802));
    outputs(668) <= layer2_outputs(4462);
    outputs(669) <= layer2_outputs(2566);
    outputs(670) <= (layer2_outputs(9247)) and not (layer2_outputs(6905));
    outputs(671) <= layer2_outputs(2295);
    outputs(672) <= layer2_outputs(8266);
    outputs(673) <= (layer2_outputs(9999)) xor (layer2_outputs(807));
    outputs(674) <= layer2_outputs(5840);
    outputs(675) <= not((layer2_outputs(4501)) and (layer2_outputs(9294)));
    outputs(676) <= layer2_outputs(4261);
    outputs(677) <= layer2_outputs(6638);
    outputs(678) <= layer2_outputs(3022);
    outputs(679) <= not(layer2_outputs(1874));
    outputs(680) <= not((layer2_outputs(6262)) xor (layer2_outputs(8099)));
    outputs(681) <= not(layer2_outputs(10012)) or (layer2_outputs(8650));
    outputs(682) <= not(layer2_outputs(4503));
    outputs(683) <= not(layer2_outputs(7285)) or (layer2_outputs(3474));
    outputs(684) <= layer2_outputs(3106);
    outputs(685) <= layer2_outputs(9046);
    outputs(686) <= not((layer2_outputs(7695)) xor (layer2_outputs(5534)));
    outputs(687) <= not(layer2_outputs(2204)) or (layer2_outputs(6604));
    outputs(688) <= layer2_outputs(1774);
    outputs(689) <= not((layer2_outputs(7138)) and (layer2_outputs(3256)));
    outputs(690) <= not(layer2_outputs(174));
    outputs(691) <= not((layer2_outputs(6902)) xor (layer2_outputs(4055)));
    outputs(692) <= not(layer2_outputs(2302));
    outputs(693) <= layer2_outputs(3937);
    outputs(694) <= layer2_outputs(9056);
    outputs(695) <= not(layer2_outputs(6941));
    outputs(696) <= not(layer2_outputs(679));
    outputs(697) <= not((layer2_outputs(8325)) xor (layer2_outputs(9795)));
    outputs(698) <= not(layer2_outputs(4302));
    outputs(699) <= layer2_outputs(2944);
    outputs(700) <= layer2_outputs(6681);
    outputs(701) <= layer2_outputs(2696);
    outputs(702) <= (layer2_outputs(7344)) xor (layer2_outputs(10065));
    outputs(703) <= (layer2_outputs(8318)) and not (layer2_outputs(715));
    outputs(704) <= layer2_outputs(5517);
    outputs(705) <= (layer2_outputs(6456)) xor (layer2_outputs(713));
    outputs(706) <= layer2_outputs(675);
    outputs(707) <= layer2_outputs(8671);
    outputs(708) <= layer2_outputs(113);
    outputs(709) <= not((layer2_outputs(7301)) or (layer2_outputs(5133)));
    outputs(710) <= (layer2_outputs(3539)) and not (layer2_outputs(6698));
    outputs(711) <= not(layer2_outputs(7789));
    outputs(712) <= not(layer2_outputs(8174));
    outputs(713) <= not((layer2_outputs(320)) xor (layer2_outputs(94)));
    outputs(714) <= (layer2_outputs(10157)) and not (layer2_outputs(647));
    outputs(715) <= not(layer2_outputs(2864));
    outputs(716) <= layer2_outputs(528);
    outputs(717) <= (layer2_outputs(5367)) and not (layer2_outputs(5587));
    outputs(718) <= (layer2_outputs(1495)) and (layer2_outputs(8472));
    outputs(719) <= not(layer2_outputs(7653));
    outputs(720) <= not(layer2_outputs(4638));
    outputs(721) <= (layer2_outputs(8337)) and (layer2_outputs(6075));
    outputs(722) <= layer2_outputs(9601);
    outputs(723) <= not(layer2_outputs(6580));
    outputs(724) <= not(layer2_outputs(4121));
    outputs(725) <= layer2_outputs(734);
    outputs(726) <= layer2_outputs(4068);
    outputs(727) <= layer2_outputs(2710);
    outputs(728) <= layer2_outputs(5548);
    outputs(729) <= not(layer2_outputs(4393));
    outputs(730) <= not(layer2_outputs(4256)) or (layer2_outputs(8506));
    outputs(731) <= layer2_outputs(4254);
    outputs(732) <= layer2_outputs(9977);
    outputs(733) <= not(layer2_outputs(9488));
    outputs(734) <= not(layer2_outputs(390));
    outputs(735) <= not(layer2_outputs(8910));
    outputs(736) <= (layer2_outputs(2380)) xor (layer2_outputs(6885));
    outputs(737) <= layer2_outputs(6881);
    outputs(738) <= not((layer2_outputs(5753)) xor (layer2_outputs(2769)));
    outputs(739) <= not(layer2_outputs(4720));
    outputs(740) <= layer2_outputs(5579);
    outputs(741) <= not(layer2_outputs(4806)) or (layer2_outputs(4826));
    outputs(742) <= (layer2_outputs(783)) and not (layer2_outputs(9821));
    outputs(743) <= (layer2_outputs(2396)) and (layer2_outputs(4356));
    outputs(744) <= not(layer2_outputs(4010));
    outputs(745) <= not(layer2_outputs(9180));
    outputs(746) <= not((layer2_outputs(4922)) xor (layer2_outputs(1287)));
    outputs(747) <= layer2_outputs(582);
    outputs(748) <= (layer2_outputs(8861)) xor (layer2_outputs(6442));
    outputs(749) <= (layer2_outputs(3443)) xor (layer2_outputs(79));
    outputs(750) <= (layer2_outputs(5367)) and not (layer2_outputs(486));
    outputs(751) <= layer2_outputs(5810);
    outputs(752) <= not(layer2_outputs(6077));
    outputs(753) <= not((layer2_outputs(8947)) xor (layer2_outputs(4237)));
    outputs(754) <= layer2_outputs(7503);
    outputs(755) <= not(layer2_outputs(5533)) or (layer2_outputs(8079));
    outputs(756) <= not(layer2_outputs(1148));
    outputs(757) <= not(layer2_outputs(4910));
    outputs(758) <= layer2_outputs(5804);
    outputs(759) <= layer2_outputs(2214);
    outputs(760) <= not(layer2_outputs(1590));
    outputs(761) <= layer2_outputs(4194);
    outputs(762) <= layer2_outputs(9895);
    outputs(763) <= layer2_outputs(5934);
    outputs(764) <= (layer2_outputs(7953)) and (layer2_outputs(9228));
    outputs(765) <= not(layer2_outputs(1639));
    outputs(766) <= not(layer2_outputs(3733)) or (layer2_outputs(3846));
    outputs(767) <= not(layer2_outputs(6565));
    outputs(768) <= not(layer2_outputs(1701));
    outputs(769) <= not((layer2_outputs(2759)) or (layer2_outputs(1308)));
    outputs(770) <= not((layer2_outputs(6400)) and (layer2_outputs(8486)));
    outputs(771) <= layer2_outputs(5596);
    outputs(772) <= (layer2_outputs(6823)) xor (layer2_outputs(8482));
    outputs(773) <= not(layer2_outputs(8351));
    outputs(774) <= layer2_outputs(7850);
    outputs(775) <= (layer2_outputs(2505)) xor (layer2_outputs(8131));
    outputs(776) <= not(layer2_outputs(3949));
    outputs(777) <= not(layer2_outputs(10069));
    outputs(778) <= layer2_outputs(5792);
    outputs(779) <= layer2_outputs(8218);
    outputs(780) <= not(layer2_outputs(9641));
    outputs(781) <= (layer2_outputs(9531)) and not (layer2_outputs(6788));
    outputs(782) <= not(layer2_outputs(1705));
    outputs(783) <= layer2_outputs(3003);
    outputs(784) <= not((layer2_outputs(6837)) xor (layer2_outputs(3364)));
    outputs(785) <= layer2_outputs(8088);
    outputs(786) <= not(layer2_outputs(8926));
    outputs(787) <= '0';
    outputs(788) <= layer2_outputs(2024);
    outputs(789) <= layer2_outputs(7647);
    outputs(790) <= not(layer2_outputs(9512));
    outputs(791) <= not(layer2_outputs(3012));
    outputs(792) <= layer2_outputs(9116);
    outputs(793) <= (layer2_outputs(3318)) and not (layer2_outputs(1885));
    outputs(794) <= not(layer2_outputs(1011));
    outputs(795) <= (layer2_outputs(1102)) and (layer2_outputs(2778));
    outputs(796) <= layer2_outputs(5472);
    outputs(797) <= (layer2_outputs(5783)) xor (layer2_outputs(969));
    outputs(798) <= not(layer2_outputs(10153));
    outputs(799) <= (layer2_outputs(5690)) xor (layer2_outputs(6216));
    outputs(800) <= not((layer2_outputs(7169)) or (layer2_outputs(5397)));
    outputs(801) <= not(layer2_outputs(3163)) or (layer2_outputs(3512));
    outputs(802) <= not((layer2_outputs(5960)) xor (layer2_outputs(9161)));
    outputs(803) <= not((layer2_outputs(9849)) xor (layer2_outputs(721)));
    outputs(804) <= not(layer2_outputs(9652));
    outputs(805) <= not(layer2_outputs(1061));
    outputs(806) <= (layer2_outputs(5781)) xor (layer2_outputs(1345));
    outputs(807) <= not(layer2_outputs(5215));
    outputs(808) <= (layer2_outputs(7798)) xor (layer2_outputs(2158));
    outputs(809) <= layer2_outputs(2421);
    outputs(810) <= (layer2_outputs(463)) xor (layer2_outputs(824));
    outputs(811) <= layer2_outputs(7595);
    outputs(812) <= not(layer2_outputs(3574));
    outputs(813) <= layer2_outputs(9713);
    outputs(814) <= (layer2_outputs(8067)) and not (layer2_outputs(3569));
    outputs(815) <= (layer2_outputs(7774)) xor (layer2_outputs(5725));
    outputs(816) <= not(layer2_outputs(4615));
    outputs(817) <= not((layer2_outputs(1986)) or (layer2_outputs(6284)));
    outputs(818) <= not(layer2_outputs(1619));
    outputs(819) <= not((layer2_outputs(1048)) xor (layer2_outputs(7230)));
    outputs(820) <= not((layer2_outputs(10020)) and (layer2_outputs(2189)));
    outputs(821) <= not(layer2_outputs(2780));
    outputs(822) <= not((layer2_outputs(8648)) or (layer2_outputs(5839)));
    outputs(823) <= not(layer2_outputs(771));
    outputs(824) <= not((layer2_outputs(6393)) xor (layer2_outputs(4373)));
    outputs(825) <= layer2_outputs(363);
    outputs(826) <= layer2_outputs(90);
    outputs(827) <= not(layer2_outputs(2706));
    outputs(828) <= not(layer2_outputs(2483));
    outputs(829) <= not((layer2_outputs(9730)) xor (layer2_outputs(3455)));
    outputs(830) <= layer2_outputs(4695);
    outputs(831) <= layer2_outputs(3449);
    outputs(832) <= (layer2_outputs(1625)) xor (layer2_outputs(8840));
    outputs(833) <= not(layer2_outputs(9677));
    outputs(834) <= not(layer2_outputs(9320));
    outputs(835) <= not((layer2_outputs(1187)) xor (layer2_outputs(1241)));
    outputs(836) <= (layer2_outputs(9946)) and (layer2_outputs(6348));
    outputs(837) <= not(layer2_outputs(8120)) or (layer2_outputs(1425));
    outputs(838) <= not(layer2_outputs(8754));
    outputs(839) <= not(layer2_outputs(9861));
    outputs(840) <= not((layer2_outputs(6241)) xor (layer2_outputs(4238)));
    outputs(841) <= layer2_outputs(1363);
    outputs(842) <= layer2_outputs(3567);
    outputs(843) <= (layer2_outputs(7422)) xor (layer2_outputs(8809));
    outputs(844) <= not(layer2_outputs(4025));
    outputs(845) <= not(layer2_outputs(7274));
    outputs(846) <= layer2_outputs(4500);
    outputs(847) <= layer2_outputs(8330);
    outputs(848) <= layer2_outputs(8906);
    outputs(849) <= not(layer2_outputs(981)) or (layer2_outputs(7148));
    outputs(850) <= not(layer2_outputs(8935));
    outputs(851) <= not((layer2_outputs(10222)) xor (layer2_outputs(9413)));
    outputs(852) <= layer2_outputs(7646);
    outputs(853) <= not((layer2_outputs(1058)) xor (layer2_outputs(8775)));
    outputs(854) <= (layer2_outputs(794)) and not (layer2_outputs(1557));
    outputs(855) <= not((layer2_outputs(1513)) xor (layer2_outputs(6855)));
    outputs(856) <= layer2_outputs(9346);
    outputs(857) <= layer2_outputs(4746);
    outputs(858) <= not(layer2_outputs(5480));
    outputs(859) <= layer2_outputs(1612);
    outputs(860) <= not(layer2_outputs(8489));
    outputs(861) <= not(layer2_outputs(2280));
    outputs(862) <= (layer2_outputs(4197)) or (layer2_outputs(7431));
    outputs(863) <= not(layer2_outputs(4259));
    outputs(864) <= not(layer2_outputs(5453)) or (layer2_outputs(9327));
    outputs(865) <= not(layer2_outputs(414));
    outputs(866) <= not(layer2_outputs(4614));
    outputs(867) <= not((layer2_outputs(2818)) xor (layer2_outputs(4486)));
    outputs(868) <= not(layer2_outputs(1380));
    outputs(869) <= layer2_outputs(1993);
    outputs(870) <= not((layer2_outputs(8054)) xor (layer2_outputs(8556)));
    outputs(871) <= not(layer2_outputs(3878));
    outputs(872) <= layer2_outputs(9772);
    outputs(873) <= (layer2_outputs(188)) xor (layer2_outputs(1575));
    outputs(874) <= not(layer2_outputs(5369));
    outputs(875) <= layer2_outputs(6172);
    outputs(876) <= layer2_outputs(7702);
    outputs(877) <= (layer2_outputs(6089)) xor (layer2_outputs(2961));
    outputs(878) <= (layer2_outputs(6816)) xor (layer2_outputs(4155));
    outputs(879) <= not((layer2_outputs(3765)) xor (layer2_outputs(3299)));
    outputs(880) <= (layer2_outputs(7737)) xor (layer2_outputs(8841));
    outputs(881) <= not((layer2_outputs(5562)) or (layer2_outputs(197)));
    outputs(882) <= not(layer2_outputs(2243));
    outputs(883) <= (layer2_outputs(62)) and not (layer2_outputs(861));
    outputs(884) <= layer2_outputs(220);
    outputs(885) <= (layer2_outputs(2676)) or (layer2_outputs(9057));
    outputs(886) <= not(layer2_outputs(2711));
    outputs(887) <= not((layer2_outputs(7247)) xor (layer2_outputs(9576)));
    outputs(888) <= (layer2_outputs(2509)) xor (layer2_outputs(8595));
    outputs(889) <= layer2_outputs(2043);
    outputs(890) <= not((layer2_outputs(1783)) xor (layer2_outputs(9079)));
    outputs(891) <= (layer2_outputs(6356)) xor (layer2_outputs(1142));
    outputs(892) <= layer2_outputs(5189);
    outputs(893) <= not(layer2_outputs(1479));
    outputs(894) <= not((layer2_outputs(5332)) or (layer2_outputs(5436)));
    outputs(895) <= not(layer2_outputs(5841));
    outputs(896) <= layer2_outputs(6715);
    outputs(897) <= not(layer2_outputs(9413)) or (layer2_outputs(7595));
    outputs(898) <= (layer2_outputs(5804)) and not (layer2_outputs(1250));
    outputs(899) <= not((layer2_outputs(1800)) and (layer2_outputs(4145)));
    outputs(900) <= not(layer2_outputs(2618));
    outputs(901) <= layer2_outputs(1507);
    outputs(902) <= not(layer2_outputs(8265));
    outputs(903) <= not(layer2_outputs(8363));
    outputs(904) <= layer2_outputs(3336);
    outputs(905) <= not((layer2_outputs(213)) xor (layer2_outputs(6315)));
    outputs(906) <= not(layer2_outputs(4220));
    outputs(907) <= not((layer2_outputs(8243)) xor (layer2_outputs(8471)));
    outputs(908) <= layer2_outputs(8191);
    outputs(909) <= not(layer2_outputs(4054)) or (layer2_outputs(1321));
    outputs(910) <= not(layer2_outputs(6774));
    outputs(911) <= layer2_outputs(2976);
    outputs(912) <= not((layer2_outputs(8317)) xor (layer2_outputs(1302)));
    outputs(913) <= layer2_outputs(10119);
    outputs(914) <= not((layer2_outputs(1058)) xor (layer2_outputs(8619)));
    outputs(915) <= layer2_outputs(817);
    outputs(916) <= layer2_outputs(336);
    outputs(917) <= layer2_outputs(8891);
    outputs(918) <= not(layer2_outputs(3140));
    outputs(919) <= layer2_outputs(8084);
    outputs(920) <= layer2_outputs(9523);
    outputs(921) <= layer2_outputs(3879);
    outputs(922) <= (layer2_outputs(2306)) xor (layer2_outputs(7245));
    outputs(923) <= layer2_outputs(2428);
    outputs(924) <= layer2_outputs(10029);
    outputs(925) <= layer2_outputs(8823);
    outputs(926) <= layer2_outputs(9552);
    outputs(927) <= not((layer2_outputs(6180)) xor (layer2_outputs(2126)));
    outputs(928) <= not(layer2_outputs(2203)) or (layer2_outputs(3653));
    outputs(929) <= not((layer2_outputs(6953)) or (layer2_outputs(7165)));
    outputs(930) <= not((layer2_outputs(7093)) xor (layer2_outputs(6639)));
    outputs(931) <= not(layer2_outputs(9927));
    outputs(932) <= not((layer2_outputs(5150)) xor (layer2_outputs(9299)));
    outputs(933) <= not(layer2_outputs(4841));
    outputs(934) <= not(layer2_outputs(2108));
    outputs(935) <= layer2_outputs(2345);
    outputs(936) <= layer2_outputs(4507);
    outputs(937) <= not(layer2_outputs(1247));
    outputs(938) <= not(layer2_outputs(286));
    outputs(939) <= not(layer2_outputs(2311)) or (layer2_outputs(3845));
    outputs(940) <= not(layer2_outputs(863));
    outputs(941) <= (layer2_outputs(8490)) xor (layer2_outputs(6874));
    outputs(942) <= layer2_outputs(479);
    outputs(943) <= not(layer2_outputs(7266));
    outputs(944) <= layer2_outputs(9272);
    outputs(945) <= not(layer2_outputs(9421));
    outputs(946) <= (layer2_outputs(6963)) and not (layer2_outputs(1498));
    outputs(947) <= not(layer2_outputs(4344));
    outputs(948) <= not(layer2_outputs(7914));
    outputs(949) <= not((layer2_outputs(626)) and (layer2_outputs(7286)));
    outputs(950) <= not(layer2_outputs(8983)) or (layer2_outputs(7732));
    outputs(951) <= not(layer2_outputs(2276)) or (layer2_outputs(9451));
    outputs(952) <= layer2_outputs(7305);
    outputs(953) <= layer2_outputs(9392);
    outputs(954) <= not(layer2_outputs(9383));
    outputs(955) <= not(layer2_outputs(10170));
    outputs(956) <= (layer2_outputs(2888)) xor (layer2_outputs(8377));
    outputs(957) <= (layer2_outputs(5265)) and not (layer2_outputs(1715));
    outputs(958) <= layer2_outputs(8700);
    outputs(959) <= layer2_outputs(1562);
    outputs(960) <= (layer2_outputs(8087)) or (layer2_outputs(9894));
    outputs(961) <= not(layer2_outputs(8951));
    outputs(962) <= (layer2_outputs(2295)) and not (layer2_outputs(2961));
    outputs(963) <= layer2_outputs(3161);
    outputs(964) <= layer2_outputs(10209);
    outputs(965) <= (layer2_outputs(6418)) and not (layer2_outputs(754));
    outputs(966) <= layer2_outputs(10171);
    outputs(967) <= (layer2_outputs(8435)) xor (layer2_outputs(2185));
    outputs(968) <= (layer2_outputs(4331)) and not (layer2_outputs(2858));
    outputs(969) <= not(layer2_outputs(4554));
    outputs(970) <= layer2_outputs(84);
    outputs(971) <= layer2_outputs(2627);
    outputs(972) <= not(layer2_outputs(5657));
    outputs(973) <= not(layer2_outputs(3360));
    outputs(974) <= (layer2_outputs(6460)) and not (layer2_outputs(9149));
    outputs(975) <= layer2_outputs(1160);
    outputs(976) <= not(layer2_outputs(8476));
    outputs(977) <= (layer2_outputs(8142)) xor (layer2_outputs(2982));
    outputs(978) <= layer2_outputs(10111);
    outputs(979) <= not(layer2_outputs(2104));
    outputs(980) <= not(layer2_outputs(573));
    outputs(981) <= (layer2_outputs(1119)) xor (layer2_outputs(9138));
    outputs(982) <= not(layer2_outputs(3249));
    outputs(983) <= (layer2_outputs(7628)) and not (layer2_outputs(4139));
    outputs(984) <= (layer2_outputs(8493)) and (layer2_outputs(4588));
    outputs(985) <= layer2_outputs(2991);
    outputs(986) <= layer2_outputs(5476);
    outputs(987) <= (layer2_outputs(10231)) and (layer2_outputs(8491));
    outputs(988) <= layer2_outputs(3562);
    outputs(989) <= not(layer2_outputs(577));
    outputs(990) <= layer2_outputs(1231);
    outputs(991) <= layer2_outputs(8742);
    outputs(992) <= not(layer2_outputs(2744));
    outputs(993) <= not(layer2_outputs(10122));
    outputs(994) <= not(layer2_outputs(1004));
    outputs(995) <= not(layer2_outputs(3260)) or (layer2_outputs(6425));
    outputs(996) <= not(layer2_outputs(116));
    outputs(997) <= not(layer2_outputs(4441));
    outputs(998) <= not(layer2_outputs(1858));
    outputs(999) <= layer2_outputs(5348);
    outputs(1000) <= (layer2_outputs(1580)) xor (layer2_outputs(2804));
    outputs(1001) <= not(layer2_outputs(9501));
    outputs(1002) <= not((layer2_outputs(2990)) xor (layer2_outputs(3893)));
    outputs(1003) <= not(layer2_outputs(10047));
    outputs(1004) <= layer2_outputs(4468);
    outputs(1005) <= layer2_outputs(8169);
    outputs(1006) <= layer2_outputs(7281);
    outputs(1007) <= not(layer2_outputs(2546));
    outputs(1008) <= not((layer2_outputs(10092)) or (layer2_outputs(8544)));
    outputs(1009) <= not(layer2_outputs(6266));
    outputs(1010) <= not(layer2_outputs(9760));
    outputs(1011) <= not(layer2_outputs(7852));
    outputs(1012) <= (layer2_outputs(433)) and (layer2_outputs(2450));
    outputs(1013) <= layer2_outputs(10105);
    outputs(1014) <= layer2_outputs(8336);
    outputs(1015) <= not(layer2_outputs(9065));
    outputs(1016) <= (layer2_outputs(10107)) xor (layer2_outputs(1189));
    outputs(1017) <= not(layer2_outputs(306));
    outputs(1018) <= (layer2_outputs(352)) and not (layer2_outputs(418));
    outputs(1019) <= not(layer2_outputs(281));
    outputs(1020) <= not((layer2_outputs(3433)) xor (layer2_outputs(9779)));
    outputs(1021) <= layer2_outputs(2777);
    outputs(1022) <= not((layer2_outputs(8123)) or (layer2_outputs(3638)));
    outputs(1023) <= not(layer2_outputs(8771)) or (layer2_outputs(5900));
    outputs(1024) <= (layer2_outputs(6721)) xor (layer2_outputs(2010));
    outputs(1025) <= not(layer2_outputs(3407));
    outputs(1026) <= not(layer2_outputs(4045));
    outputs(1027) <= layer2_outputs(5234);
    outputs(1028) <= not(layer2_outputs(1235));
    outputs(1029) <= not((layer2_outputs(4368)) xor (layer2_outputs(109)));
    outputs(1030) <= not((layer2_outputs(3517)) xor (layer2_outputs(6864)));
    outputs(1031) <= not(layer2_outputs(8673));
    outputs(1032) <= not(layer2_outputs(5741));
    outputs(1033) <= (layer2_outputs(7485)) and not (layer2_outputs(4954));
    outputs(1034) <= layer2_outputs(3316);
    outputs(1035) <= not(layer2_outputs(6879));
    outputs(1036) <= not((layer2_outputs(3129)) xor (layer2_outputs(7307)));
    outputs(1037) <= not(layer2_outputs(10146));
    outputs(1038) <= layer2_outputs(5394);
    outputs(1039) <= (layer2_outputs(482)) and (layer2_outputs(9114));
    outputs(1040) <= (layer2_outputs(8507)) and not (layer2_outputs(8051));
    outputs(1041) <= (layer2_outputs(1211)) xor (layer2_outputs(1188));
    outputs(1042) <= not((layer2_outputs(4589)) xor (layer2_outputs(8207)));
    outputs(1043) <= (layer2_outputs(9034)) xor (layer2_outputs(5152));
    outputs(1044) <= not(layer2_outputs(3005));
    outputs(1045) <= not(layer2_outputs(8248));
    outputs(1046) <= not(layer2_outputs(5488));
    outputs(1047) <= not((layer2_outputs(8627)) or (layer2_outputs(9384)));
    outputs(1048) <= (layer2_outputs(3178)) and not (layer2_outputs(2116));
    outputs(1049) <= (layer2_outputs(3079)) and not (layer2_outputs(2717));
    outputs(1050) <= not((layer2_outputs(5912)) or (layer2_outputs(342)));
    outputs(1051) <= (layer2_outputs(3704)) or (layer2_outputs(9242));
    outputs(1052) <= layer2_outputs(1037);
    outputs(1053) <= (layer2_outputs(10119)) xor (layer2_outputs(7821));
    outputs(1054) <= (layer2_outputs(5799)) and not (layer2_outputs(6012));
    outputs(1055) <= (layer2_outputs(4729)) and not (layer2_outputs(7702));
    outputs(1056) <= (layer2_outputs(6772)) and (layer2_outputs(6511));
    outputs(1057) <= not(layer2_outputs(7076)) or (layer2_outputs(9452));
    outputs(1058) <= not((layer2_outputs(2752)) or (layer2_outputs(5877)));
    outputs(1059) <= (layer2_outputs(3812)) xor (layer2_outputs(842));
    outputs(1060) <= not(layer2_outputs(3587));
    outputs(1061) <= not((layer2_outputs(6451)) xor (layer2_outputs(5951)));
    outputs(1062) <= not((layer2_outputs(4926)) or (layer2_outputs(6708)));
    outputs(1063) <= not((layer2_outputs(10011)) xor (layer2_outputs(10204)));
    outputs(1064) <= (layer2_outputs(7125)) xor (layer2_outputs(9685));
    outputs(1065) <= not(layer2_outputs(5831));
    outputs(1066) <= (layer2_outputs(1577)) xor (layer2_outputs(7211));
    outputs(1067) <= (layer2_outputs(6562)) xor (layer2_outputs(9687));
    outputs(1068) <= (layer2_outputs(7040)) xor (layer2_outputs(4744));
    outputs(1069) <= (layer2_outputs(707)) xor (layer2_outputs(9980));
    outputs(1070) <= (layer2_outputs(8100)) and not (layer2_outputs(7399));
    outputs(1071) <= (layer2_outputs(7944)) and not (layer2_outputs(4107));
    outputs(1072) <= (layer2_outputs(8770)) xor (layer2_outputs(9899));
    outputs(1073) <= not((layer2_outputs(3148)) xor (layer2_outputs(5756)));
    outputs(1074) <= (layer2_outputs(5386)) or (layer2_outputs(7343));
    outputs(1075) <= layer2_outputs(6245);
    outputs(1076) <= layer2_outputs(7057);
    outputs(1077) <= not(layer2_outputs(9575));
    outputs(1078) <= (layer2_outputs(9000)) and not (layer2_outputs(8234));
    outputs(1079) <= (layer2_outputs(8744)) and (layer2_outputs(631));
    outputs(1080) <= (layer2_outputs(3582)) and not (layer2_outputs(2292));
    outputs(1081) <= (layer2_outputs(3131)) and not (layer2_outputs(6274));
    outputs(1082) <= layer2_outputs(3206);
    outputs(1083) <= (layer2_outputs(8437)) and (layer2_outputs(9318));
    outputs(1084) <= (layer2_outputs(7407)) and not (layer2_outputs(8588));
    outputs(1085) <= not((layer2_outputs(1089)) xor (layer2_outputs(7522)));
    outputs(1086) <= not((layer2_outputs(7518)) or (layer2_outputs(7268)));
    outputs(1087) <= layer2_outputs(6533);
    outputs(1088) <= not(layer2_outputs(2824));
    outputs(1089) <= not((layer2_outputs(9604)) xor (layer2_outputs(6211)));
    outputs(1090) <= (layer2_outputs(4500)) xor (layer2_outputs(2644));
    outputs(1091) <= (layer2_outputs(9907)) xor (layer2_outputs(3592));
    outputs(1092) <= not((layer2_outputs(5121)) xor (layer2_outputs(7624)));
    outputs(1093) <= not((layer2_outputs(950)) or (layer2_outputs(433)));
    outputs(1094) <= (layer2_outputs(1228)) xor (layer2_outputs(8395));
    outputs(1095) <= (layer2_outputs(9891)) and (layer2_outputs(5157));
    outputs(1096) <= not((layer2_outputs(9938)) or (layer2_outputs(8929)));
    outputs(1097) <= (layer2_outputs(9661)) xor (layer2_outputs(4860));
    outputs(1098) <= '0';
    outputs(1099) <= not(layer2_outputs(2267));
    outputs(1100) <= not(layer2_outputs(5017));
    outputs(1101) <= (layer2_outputs(9416)) and (layer2_outputs(210));
    outputs(1102) <= not(layer2_outputs(9243));
    outputs(1103) <= not(layer2_outputs(10145));
    outputs(1104) <= (layer2_outputs(2393)) xor (layer2_outputs(2206));
    outputs(1105) <= layer2_outputs(5477);
    outputs(1106) <= not((layer2_outputs(8150)) or (layer2_outputs(5913)));
    outputs(1107) <= layer2_outputs(2171);
    outputs(1108) <= (layer2_outputs(2176)) and (layer2_outputs(5303));
    outputs(1109) <= not((layer2_outputs(5914)) xor (layer2_outputs(2403)));
    outputs(1110) <= (layer2_outputs(1011)) and (layer2_outputs(1629));
    outputs(1111) <= (layer2_outputs(282)) and not (layer2_outputs(4509));
    outputs(1112) <= not((layer2_outputs(6575)) or (layer2_outputs(2861)));
    outputs(1113) <= (layer2_outputs(7135)) and (layer2_outputs(2384));
    outputs(1114) <= not(layer2_outputs(8283));
    outputs(1115) <= layer2_outputs(2177);
    outputs(1116) <= (layer2_outputs(9535)) xor (layer2_outputs(7968));
    outputs(1117) <= (layer2_outputs(6485)) xor (layer2_outputs(7616));
    outputs(1118) <= not(layer2_outputs(4988));
    outputs(1119) <= (layer2_outputs(8497)) and (layer2_outputs(2071));
    outputs(1120) <= layer2_outputs(8214);
    outputs(1121) <= (layer2_outputs(4395)) xor (layer2_outputs(4829));
    outputs(1122) <= (layer2_outputs(6756)) and not (layer2_outputs(9108));
    outputs(1123) <= layer2_outputs(3483);
    outputs(1124) <= not((layer2_outputs(8435)) xor (layer2_outputs(905)));
    outputs(1125) <= layer2_outputs(5328);
    outputs(1126) <= (layer2_outputs(746)) xor (layer2_outputs(7747));
    outputs(1127) <= not(layer2_outputs(8133));
    outputs(1128) <= not(layer2_outputs(3561));
    outputs(1129) <= not(layer2_outputs(2514));
    outputs(1130) <= not((layer2_outputs(8610)) xor (layer2_outputs(5441)));
    outputs(1131) <= layer2_outputs(1290);
    outputs(1132) <= layer2_outputs(4891);
    outputs(1133) <= layer2_outputs(9173);
    outputs(1134) <= not((layer2_outputs(1238)) xor (layer2_outputs(2893)));
    outputs(1135) <= layer2_outputs(326);
    outputs(1136) <= not((layer2_outputs(3066)) or (layer2_outputs(672)));
    outputs(1137) <= layer2_outputs(2709);
    outputs(1138) <= layer2_outputs(87);
    outputs(1139) <= layer2_outputs(6219);
    outputs(1140) <= layer2_outputs(9993);
    outputs(1141) <= (layer2_outputs(7332)) xor (layer2_outputs(5359));
    outputs(1142) <= not(layer2_outputs(1770));
    outputs(1143) <= (layer2_outputs(87)) and not (layer2_outputs(2996));
    outputs(1144) <= not((layer2_outputs(9243)) xor (layer2_outputs(2889)));
    outputs(1145) <= (layer2_outputs(6359)) xor (layer2_outputs(8017));
    outputs(1146) <= layer2_outputs(2115);
    outputs(1147) <= not(layer2_outputs(9704));
    outputs(1148) <= not(layer2_outputs(3597));
    outputs(1149) <= not((layer2_outputs(3913)) xor (layer2_outputs(651)));
    outputs(1150) <= layer2_outputs(347);
    outputs(1151) <= layer2_outputs(4850);
    outputs(1152) <= not((layer2_outputs(3429)) or (layer2_outputs(10021)));
    outputs(1153) <= layer2_outputs(5080);
    outputs(1154) <= not(layer2_outputs(3384));
    outputs(1155) <= not((layer2_outputs(520)) xor (layer2_outputs(1223)));
    outputs(1156) <= layer2_outputs(5946);
    outputs(1157) <= not(layer2_outputs(10093)) or (layer2_outputs(2014));
    outputs(1158) <= not((layer2_outputs(1460)) xor (layer2_outputs(2716)));
    outputs(1159) <= layer2_outputs(4609);
    outputs(1160) <= (layer2_outputs(8816)) and (layer2_outputs(6102));
    outputs(1161) <= (layer2_outputs(429)) xor (layer2_outputs(2760));
    outputs(1162) <= (layer2_outputs(7711)) and not (layer2_outputs(4534));
    outputs(1163) <= not((layer2_outputs(10159)) xor (layer2_outputs(5924)));
    outputs(1164) <= not(layer2_outputs(7935));
    outputs(1165) <= (layer2_outputs(2066)) and not (layer2_outputs(9745));
    outputs(1166) <= layer2_outputs(1010);
    outputs(1167) <= not((layer2_outputs(5615)) xor (layer2_outputs(5532)));
    outputs(1168) <= not(layer2_outputs(4455));
    outputs(1169) <= (layer2_outputs(4775)) xor (layer2_outputs(9216));
    outputs(1170) <= (layer2_outputs(5812)) and (layer2_outputs(6218));
    outputs(1171) <= layer2_outputs(593);
    outputs(1172) <= not(layer2_outputs(5821));
    outputs(1173) <= (layer2_outputs(4664)) and (layer2_outputs(3776));
    outputs(1174) <= not(layer2_outputs(10031));
    outputs(1175) <= layer2_outputs(8560);
    outputs(1176) <= (layer2_outputs(1945)) and not (layer2_outputs(8548));
    outputs(1177) <= layer2_outputs(476);
    outputs(1178) <= (layer2_outputs(5144)) xor (layer2_outputs(9787));
    outputs(1179) <= (layer2_outputs(6143)) and (layer2_outputs(755));
    outputs(1180) <= (layer2_outputs(283)) and (layer2_outputs(5897));
    outputs(1181) <= (layer2_outputs(973)) and (layer2_outputs(10208));
    outputs(1182) <= layer2_outputs(7154);
    outputs(1183) <= not(layer2_outputs(5922));
    outputs(1184) <= layer2_outputs(2920);
    outputs(1185) <= not(layer2_outputs(1482));
    outputs(1186) <= layer2_outputs(1692);
    outputs(1187) <= (layer2_outputs(9183)) or (layer2_outputs(2829));
    outputs(1188) <= (layer2_outputs(7406)) and (layer2_outputs(1954));
    outputs(1189) <= (layer2_outputs(6480)) and (layer2_outputs(10136));
    outputs(1190) <= not((layer2_outputs(5714)) xor (layer2_outputs(9929)));
    outputs(1191) <= not(layer2_outputs(7078));
    outputs(1192) <= (layer2_outputs(8604)) and not (layer2_outputs(2844));
    outputs(1193) <= not((layer2_outputs(713)) or (layer2_outputs(3120)));
    outputs(1194) <= not((layer2_outputs(10228)) xor (layer2_outputs(6450)));
    outputs(1195) <= not((layer2_outputs(3851)) xor (layer2_outputs(8541)));
    outputs(1196) <= not(layer2_outputs(1781));
    outputs(1197) <= (layer2_outputs(3550)) xor (layer2_outputs(3634));
    outputs(1198) <= not((layer2_outputs(2683)) xor (layer2_outputs(8434)));
    outputs(1199) <= layer2_outputs(9017);
    outputs(1200) <= not((layer2_outputs(7474)) or (layer2_outputs(6313)));
    outputs(1201) <= not(layer2_outputs(3393));
    outputs(1202) <= not(layer2_outputs(5947));
    outputs(1203) <= not((layer2_outputs(9809)) or (layer2_outputs(7338)));
    outputs(1204) <= layer2_outputs(2125);
    outputs(1205) <= not(layer2_outputs(9474));
    outputs(1206) <= not((layer2_outputs(7381)) or (layer2_outputs(3599)));
    outputs(1207) <= not(layer2_outputs(9992));
    outputs(1208) <= (layer2_outputs(5926)) xor (layer2_outputs(762));
    outputs(1209) <= (layer2_outputs(1225)) and (layer2_outputs(235));
    outputs(1210) <= not(layer2_outputs(4239));
    outputs(1211) <= (layer2_outputs(6029)) and not (layer2_outputs(2181));
    outputs(1212) <= layer2_outputs(546);
    outputs(1213) <= (layer2_outputs(5583)) and (layer2_outputs(1835));
    outputs(1214) <= not((layer2_outputs(3383)) xor (layer2_outputs(6379)));
    outputs(1215) <= not((layer2_outputs(3218)) xor (layer2_outputs(9691)));
    outputs(1216) <= (layer2_outputs(6962)) xor (layer2_outputs(7613));
    outputs(1217) <= (layer2_outputs(7253)) and not (layer2_outputs(7205));
    outputs(1218) <= not((layer2_outputs(7682)) xor (layer2_outputs(378)));
    outputs(1219) <= layer2_outputs(4731);
    outputs(1220) <= layer2_outputs(5355);
    outputs(1221) <= not((layer2_outputs(10198)) or (layer2_outputs(7151)));
    outputs(1222) <= layer2_outputs(4233);
    outputs(1223) <= not(layer2_outputs(3390));
    outputs(1224) <= (layer2_outputs(8979)) and not (layer2_outputs(4532));
    outputs(1225) <= layer2_outputs(7241);
    outputs(1226) <= not(layer2_outputs(6253));
    outputs(1227) <= (layer2_outputs(7608)) and not (layer2_outputs(9200));
    outputs(1228) <= not(layer2_outputs(4582));
    outputs(1229) <= (layer2_outputs(3768)) xor (layer2_outputs(8694));
    outputs(1230) <= layer2_outputs(1885);
    outputs(1231) <= (layer2_outputs(1687)) and (layer2_outputs(7372));
    outputs(1232) <= not(layer2_outputs(7020));
    outputs(1233) <= layer2_outputs(3089);
    outputs(1234) <= not(layer2_outputs(6909));
    outputs(1235) <= not(layer2_outputs(5422));
    outputs(1236) <= not((layer2_outputs(3456)) or (layer2_outputs(5130)));
    outputs(1237) <= (layer2_outputs(4504)) and not (layer2_outputs(9207));
    outputs(1238) <= not(layer2_outputs(4228));
    outputs(1239) <= (layer2_outputs(3058)) and not (layer2_outputs(3508));
    outputs(1240) <= not(layer2_outputs(1680));
    outputs(1241) <= layer2_outputs(7242);
    outputs(1242) <= layer2_outputs(9041);
    outputs(1243) <= not((layer2_outputs(2219)) xor (layer2_outputs(8328)));
    outputs(1244) <= layer2_outputs(6143);
    outputs(1245) <= not(layer2_outputs(9437));
    outputs(1246) <= (layer2_outputs(1051)) xor (layer2_outputs(6066));
    outputs(1247) <= (layer2_outputs(2782)) xor (layer2_outputs(9679));
    outputs(1248) <= (layer2_outputs(2049)) and (layer2_outputs(2392));
    outputs(1249) <= not(layer2_outputs(4800));
    outputs(1250) <= layer2_outputs(2720);
    outputs(1251) <= (layer2_outputs(3748)) and (layer2_outputs(83));
    outputs(1252) <= (layer2_outputs(6121)) and (layer2_outputs(10167));
    outputs(1253) <= not(layer2_outputs(3048));
    outputs(1254) <= layer2_outputs(7166);
    outputs(1255) <= not(layer2_outputs(3840));
    outputs(1256) <= not((layer2_outputs(6306)) xor (layer2_outputs(3370)));
    outputs(1257) <= (layer2_outputs(6298)) xor (layer2_outputs(1985));
    outputs(1258) <= not((layer2_outputs(3715)) xor (layer2_outputs(4863)));
    outputs(1259) <= (layer2_outputs(3013)) and (layer2_outputs(4108));
    outputs(1260) <= (layer2_outputs(2826)) xor (layer2_outputs(4085));
    outputs(1261) <= layer2_outputs(3669);
    outputs(1262) <= layer2_outputs(4172);
    outputs(1263) <= not(layer2_outputs(3574));
    outputs(1264) <= (layer2_outputs(9686)) xor (layer2_outputs(3541));
    outputs(1265) <= layer2_outputs(2924);
    outputs(1266) <= not(layer2_outputs(7731));
    outputs(1267) <= layer2_outputs(4184);
    outputs(1268) <= not((layer2_outputs(7703)) xor (layer2_outputs(1668)));
    outputs(1269) <= layer2_outputs(5233);
    outputs(1270) <= (layer2_outputs(5727)) xor (layer2_outputs(9780));
    outputs(1271) <= (layer2_outputs(8771)) xor (layer2_outputs(9097));
    outputs(1272) <= not(layer2_outputs(7713));
    outputs(1273) <= not((layer2_outputs(2131)) xor (layer2_outputs(6656)));
    outputs(1274) <= (layer2_outputs(1625)) and not (layer2_outputs(2707));
    outputs(1275) <= (layer2_outputs(6249)) and (layer2_outputs(3139));
    outputs(1276) <= (layer2_outputs(8708)) xor (layer2_outputs(1595));
    outputs(1277) <= not(layer2_outputs(5075));
    outputs(1278) <= not(layer2_outputs(8804));
    outputs(1279) <= not((layer2_outputs(140)) xor (layer2_outputs(4444)));
    outputs(1280) <= (layer2_outputs(6539)) and (layer2_outputs(8960));
    outputs(1281) <= not((layer2_outputs(3092)) and (layer2_outputs(9152)));
    outputs(1282) <= not((layer2_outputs(8368)) xor (layer2_outputs(7988)));
    outputs(1283) <= not((layer2_outputs(7496)) xor (layer2_outputs(5739)));
    outputs(1284) <= layer2_outputs(3640);
    outputs(1285) <= (layer2_outputs(4844)) xor (layer2_outputs(6862));
    outputs(1286) <= (layer2_outputs(4306)) and not (layer2_outputs(3647));
    outputs(1287) <= (layer2_outputs(3086)) xor (layer2_outputs(8311));
    outputs(1288) <= not(layer2_outputs(2269)) or (layer2_outputs(7998));
    outputs(1289) <= not(layer2_outputs(4809));
    outputs(1290) <= not(layer2_outputs(8));
    outputs(1291) <= layer2_outputs(173);
    outputs(1292) <= not(layer2_outputs(4509));
    outputs(1293) <= (layer2_outputs(2261)) xor (layer2_outputs(2828));
    outputs(1294) <= not((layer2_outputs(3948)) and (layer2_outputs(5083)));
    outputs(1295) <= (layer2_outputs(2300)) and not (layer2_outputs(1586));
    outputs(1296) <= not(layer2_outputs(747));
    outputs(1297) <= layer2_outputs(9958);
    outputs(1298) <= not((layer2_outputs(2838)) xor (layer2_outputs(1643)));
    outputs(1299) <= not(layer2_outputs(6230));
    outputs(1300) <= (layer2_outputs(7910)) and not (layer2_outputs(4687));
    outputs(1301) <= not((layer2_outputs(4822)) xor (layer2_outputs(9644)));
    outputs(1302) <= (layer2_outputs(6946)) and not (layer2_outputs(9750));
    outputs(1303) <= (layer2_outputs(6747)) and not (layer2_outputs(5225));
    outputs(1304) <= not(layer2_outputs(1283));
    outputs(1305) <= (layer2_outputs(5920)) and (layer2_outputs(8364));
    outputs(1306) <= layer2_outputs(7666);
    outputs(1307) <= (layer2_outputs(2324)) and not (layer2_outputs(6441));
    outputs(1308) <= not(layer2_outputs(9909));
    outputs(1309) <= (layer2_outputs(6790)) xor (layer2_outputs(1415));
    outputs(1310) <= layer2_outputs(3382);
    outputs(1311) <= layer2_outputs(9369);
    outputs(1312) <= not((layer2_outputs(8289)) or (layer2_outputs(2976)));
    outputs(1313) <= not(layer2_outputs(8014)) or (layer2_outputs(5005));
    outputs(1314) <= (layer2_outputs(10188)) and not (layer2_outputs(4561));
    outputs(1315) <= (layer2_outputs(7637)) and (layer2_outputs(7163));
    outputs(1316) <= not(layer2_outputs(2473));
    outputs(1317) <= not((layer2_outputs(6849)) or (layer2_outputs(10173)));
    outputs(1318) <= layer2_outputs(1070);
    outputs(1319) <= not(layer2_outputs(5481));
    outputs(1320) <= not(layer2_outputs(9424));
    outputs(1321) <= (layer2_outputs(117)) and not (layer2_outputs(8830));
    outputs(1322) <= not((layer2_outputs(1374)) xor (layer2_outputs(8749)));
    outputs(1323) <= not((layer2_outputs(5290)) or (layer2_outputs(6038)));
    outputs(1324) <= not((layer2_outputs(3255)) xor (layer2_outputs(3227)));
    outputs(1325) <= not((layer2_outputs(1337)) or (layer2_outputs(4941)));
    outputs(1326) <= not(layer2_outputs(8205));
    outputs(1327) <= not((layer2_outputs(897)) or (layer2_outputs(9623)));
    outputs(1328) <= not(layer2_outputs(3409));
    outputs(1329) <= layer2_outputs(464);
    outputs(1330) <= not(layer2_outputs(6971));
    outputs(1331) <= not((layer2_outputs(6560)) xor (layer2_outputs(7641)));
    outputs(1332) <= (layer2_outputs(808)) xor (layer2_outputs(8515));
    outputs(1333) <= layer2_outputs(5523);
    outputs(1334) <= not((layer2_outputs(4408)) and (layer2_outputs(7715)));
    outputs(1335) <= '0';
    outputs(1336) <= not(layer2_outputs(1979));
    outputs(1337) <= layer2_outputs(3301);
    outputs(1338) <= (layer2_outputs(3589)) and not (layer2_outputs(3675));
    outputs(1339) <= layer2_outputs(9869);
    outputs(1340) <= layer2_outputs(2494);
    outputs(1341) <= (layer2_outputs(8617)) and (layer2_outputs(8599));
    outputs(1342) <= layer2_outputs(5326);
    outputs(1343) <= layer2_outputs(5239);
    outputs(1344) <= not((layer2_outputs(5090)) xor (layer2_outputs(9735)));
    outputs(1345) <= not((layer2_outputs(5528)) xor (layer2_outputs(9262)));
    outputs(1346) <= (layer2_outputs(5748)) and (layer2_outputs(8539));
    outputs(1347) <= not((layer2_outputs(8441)) xor (layer2_outputs(6992)));
    outputs(1348) <= not(layer2_outputs(4691));
    outputs(1349) <= not((layer2_outputs(5124)) and (layer2_outputs(7023)));
    outputs(1350) <= not(layer2_outputs(8837));
    outputs(1351) <= not((layer2_outputs(8198)) or (layer2_outputs(9768)));
    outputs(1352) <= layer2_outputs(5761);
    outputs(1353) <= (layer2_outputs(5058)) or (layer2_outputs(8032));
    outputs(1354) <= not((layer2_outputs(7306)) xor (layer2_outputs(8056)));
    outputs(1355) <= not(layer2_outputs(5928));
    outputs(1356) <= not(layer2_outputs(1409));
    outputs(1357) <= not(layer2_outputs(5409));
    outputs(1358) <= not((layer2_outputs(6843)) or (layer2_outputs(2248)));
    outputs(1359) <= not((layer2_outputs(1040)) xor (layer2_outputs(2722)));
    outputs(1360) <= not(layer2_outputs(7085));
    outputs(1361) <= layer2_outputs(2708);
    outputs(1362) <= layer2_outputs(3831);
    outputs(1363) <= not(layer2_outputs(5065));
    outputs(1364) <= not(layer2_outputs(2862));
    outputs(1365) <= layer2_outputs(6459);
    outputs(1366) <= layer2_outputs(1029);
    outputs(1367) <= not((layer2_outputs(4268)) xor (layer2_outputs(2349)));
    outputs(1368) <= not((layer2_outputs(7319)) or (layer2_outputs(8221)));
    outputs(1369) <= not((layer2_outputs(6683)) xor (layer2_outputs(7504)));
    outputs(1370) <= not((layer2_outputs(10065)) or (layer2_outputs(6018)));
    outputs(1371) <= layer2_outputs(5729);
    outputs(1372) <= (layer2_outputs(9690)) xor (layer2_outputs(9491));
    outputs(1373) <= not(layer2_outputs(3130));
    outputs(1374) <= not(layer2_outputs(9128));
    outputs(1375) <= (layer2_outputs(1685)) and not (layer2_outputs(214));
    outputs(1376) <= (layer2_outputs(7826)) and (layer2_outputs(5817));
    outputs(1377) <= not(layer2_outputs(300));
    outputs(1378) <= (layer2_outputs(710)) and not (layer2_outputs(3082));
    outputs(1379) <= not(layer2_outputs(1193));
    outputs(1380) <= not((layer2_outputs(7916)) or (layer2_outputs(6719)));
    outputs(1381) <= (layer2_outputs(4681)) and (layer2_outputs(4583));
    outputs(1382) <= not(layer2_outputs(5265)) or (layer2_outputs(3506));
    outputs(1383) <= (layer2_outputs(414)) xor (layer2_outputs(456));
    outputs(1384) <= not((layer2_outputs(8856)) or (layer2_outputs(9783)));
    outputs(1385) <= layer2_outputs(1023);
    outputs(1386) <= not(layer2_outputs(4539));
    outputs(1387) <= not(layer2_outputs(3680));
    outputs(1388) <= (layer2_outputs(7894)) xor (layer2_outputs(8974));
    outputs(1389) <= not(layer2_outputs(9740));
    outputs(1390) <= (layer2_outputs(8203)) and not (layer2_outputs(5177));
    outputs(1391) <= layer2_outputs(4161);
    outputs(1392) <= layer2_outputs(7068);
    outputs(1393) <= not(layer2_outputs(8269));
    outputs(1394) <= (layer2_outputs(3129)) and (layer2_outputs(6934));
    outputs(1395) <= (layer2_outputs(7047)) xor (layer2_outputs(4823));
    outputs(1396) <= not(layer2_outputs(4361));
    outputs(1397) <= (layer2_outputs(8691)) and (layer2_outputs(8244));
    outputs(1398) <= not((layer2_outputs(7281)) xor (layer2_outputs(7478)));
    outputs(1399) <= not((layer2_outputs(4492)) or (layer2_outputs(6076)));
    outputs(1400) <= (layer2_outputs(7344)) xor (layer2_outputs(6151));
    outputs(1401) <= layer2_outputs(6132);
    outputs(1402) <= not(layer2_outputs(2700));
    outputs(1403) <= not(layer2_outputs(3305));
    outputs(1404) <= not(layer2_outputs(9332));
    outputs(1405) <= not((layer2_outputs(5472)) xor (layer2_outputs(3485)));
    outputs(1406) <= (layer2_outputs(7774)) and (layer2_outputs(2763));
    outputs(1407) <= not(layer2_outputs(6307));
    outputs(1408) <= (layer2_outputs(530)) xor (layer2_outputs(9615));
    outputs(1409) <= not(layer2_outputs(8597));
    outputs(1410) <= not(layer2_outputs(8099));
    outputs(1411) <= (layer2_outputs(4515)) xor (layer2_outputs(799));
    outputs(1412) <= layer2_outputs(5723);
    outputs(1413) <= not(layer2_outputs(5048)) or (layer2_outputs(1360));
    outputs(1414) <= layer2_outputs(170);
    outputs(1415) <= (layer2_outputs(574)) or (layer2_outputs(2092));
    outputs(1416) <= (layer2_outputs(1927)) and not (layer2_outputs(5452));
    outputs(1417) <= not((layer2_outputs(5193)) xor (layer2_outputs(5970)));
    outputs(1418) <= not(layer2_outputs(3614));
    outputs(1419) <= layer2_outputs(889);
    outputs(1420) <= not((layer2_outputs(1165)) xor (layer2_outputs(4779)));
    outputs(1421) <= layer2_outputs(4494);
    outputs(1422) <= not((layer2_outputs(9746)) xor (layer2_outputs(6009)));
    outputs(1423) <= not(layer2_outputs(4873));
    outputs(1424) <= not(layer2_outputs(8133));
    outputs(1425) <= layer2_outputs(7193);
    outputs(1426) <= (layer2_outputs(7416)) and not (layer2_outputs(5709));
    outputs(1427) <= (layer2_outputs(232)) xor (layer2_outputs(6673));
    outputs(1428) <= (layer2_outputs(5919)) and (layer2_outputs(2994));
    outputs(1429) <= (layer2_outputs(9926)) xor (layer2_outputs(3136));
    outputs(1430) <= layer2_outputs(9158);
    outputs(1431) <= not(layer2_outputs(10010));
    outputs(1432) <= (layer2_outputs(9500)) and (layer2_outputs(5552));
    outputs(1433) <= (layer2_outputs(1416)) xor (layer2_outputs(6742));
    outputs(1434) <= not((layer2_outputs(3593)) xor (layer2_outputs(2336)));
    outputs(1435) <= (layer2_outputs(9290)) and not (layer2_outputs(6543));
    outputs(1436) <= (layer2_outputs(5885)) xor (layer2_outputs(888));
    outputs(1437) <= layer2_outputs(6582);
    outputs(1438) <= not(layer2_outputs(5339));
    outputs(1439) <= (layer2_outputs(7239)) and not (layer2_outputs(5955));
    outputs(1440) <= (layer2_outputs(5753)) and not (layer2_outputs(2275));
    outputs(1441) <= layer2_outputs(7143);
    outputs(1442) <= (layer2_outputs(8669)) xor (layer2_outputs(3163));
    outputs(1443) <= layer2_outputs(8008);
    outputs(1444) <= not((layer2_outputs(986)) xor (layer2_outputs(533)));
    outputs(1445) <= layer2_outputs(5860);
    outputs(1446) <= '0';
    outputs(1447) <= not((layer2_outputs(1200)) xor (layer2_outputs(3118)));
    outputs(1448) <= (layer2_outputs(9022)) and not (layer2_outputs(2139));
    outputs(1449) <= (layer2_outputs(3087)) xor (layer2_outputs(9687));
    outputs(1450) <= (layer2_outputs(6757)) and not (layer2_outputs(241));
    outputs(1451) <= (layer2_outputs(9068)) or (layer2_outputs(5309));
    outputs(1452) <= not(layer2_outputs(3727));
    outputs(1453) <= layer2_outputs(9480);
    outputs(1454) <= layer2_outputs(1343);
    outputs(1455) <= not((layer2_outputs(9190)) xor (layer2_outputs(2667)));
    outputs(1456) <= (layer2_outputs(776)) and not (layer2_outputs(1285));
    outputs(1457) <= layer2_outputs(561);
    outputs(1458) <= not(layer2_outputs(5605));
    outputs(1459) <= (layer2_outputs(6481)) xor (layer2_outputs(161));
    outputs(1460) <= not(layer2_outputs(9544));
    outputs(1461) <= not((layer2_outputs(2329)) or (layer2_outputs(10100)));
    outputs(1462) <= layer2_outputs(7779);
    outputs(1463) <= (layer2_outputs(2843)) or (layer2_outputs(1880));
    outputs(1464) <= layer2_outputs(6684);
    outputs(1465) <= not(layer2_outputs(10058)) or (layer2_outputs(2327));
    outputs(1466) <= (layer2_outputs(9017)) and not (layer2_outputs(6668));
    outputs(1467) <= (layer2_outputs(619)) and (layer2_outputs(9110));
    outputs(1468) <= (layer2_outputs(2412)) and (layer2_outputs(9910));
    outputs(1469) <= not((layer2_outputs(5045)) or (layer2_outputs(1374)));
    outputs(1470) <= (layer2_outputs(9645)) and not (layer2_outputs(7988));
    outputs(1471) <= layer2_outputs(7419);
    outputs(1472) <= not(layer2_outputs(6827));
    outputs(1473) <= not(layer2_outputs(3243));
    outputs(1474) <= not((layer2_outputs(8835)) xor (layer2_outputs(5142)));
    outputs(1475) <= not((layer2_outputs(8418)) xor (layer2_outputs(491)));
    outputs(1476) <= (layer2_outputs(6131)) and not (layer2_outputs(10132));
    outputs(1477) <= layer2_outputs(5194);
    outputs(1478) <= (layer2_outputs(5843)) and (layer2_outputs(5515));
    outputs(1479) <= not((layer2_outputs(4167)) xor (layer2_outputs(7016)));
    outputs(1480) <= (layer2_outputs(7056)) and (layer2_outputs(8746));
    outputs(1481) <= (layer2_outputs(1361)) xor (layer2_outputs(4950));
    outputs(1482) <= not(layer2_outputs(5210)) or (layer2_outputs(8510));
    outputs(1483) <= not(layer2_outputs(3991));
    outputs(1484) <= (layer2_outputs(5129)) and not (layer2_outputs(4635));
    outputs(1485) <= (layer2_outputs(8824)) xor (layer2_outputs(3507));
    outputs(1486) <= not(layer2_outputs(3409));
    outputs(1487) <= (layer2_outputs(5371)) and not (layer2_outputs(4151));
    outputs(1488) <= not(layer2_outputs(7451));
    outputs(1489) <= layer2_outputs(5289);
    outputs(1490) <= (layer2_outputs(4641)) xor (layer2_outputs(8635));
    outputs(1491) <= not((layer2_outputs(8778)) xor (layer2_outputs(6427)));
    outputs(1492) <= layer2_outputs(5490);
    outputs(1493) <= not(layer2_outputs(3254)) or (layer2_outputs(10161));
    outputs(1494) <= not((layer2_outputs(417)) xor (layer2_outputs(2766)));
    outputs(1495) <= layer2_outputs(8353);
    outputs(1496) <= not((layer2_outputs(8563)) xor (layer2_outputs(8612)));
    outputs(1497) <= layer2_outputs(1410);
    outputs(1498) <= (layer2_outputs(5609)) and (layer2_outputs(10196));
    outputs(1499) <= layer2_outputs(3421);
    outputs(1500) <= layer2_outputs(1190);
    outputs(1501) <= (layer2_outputs(6366)) xor (layer2_outputs(7851));
    outputs(1502) <= layer2_outputs(7267);
    outputs(1503) <= not(layer2_outputs(8967));
    outputs(1504) <= layer2_outputs(5200);
    outputs(1505) <= (layer2_outputs(3930)) and (layer2_outputs(5251));
    outputs(1506) <= not(layer2_outputs(7785));
    outputs(1507) <= layer2_outputs(9769);
    outputs(1508) <= not((layer2_outputs(3402)) xor (layer2_outputs(7511)));
    outputs(1509) <= not((layer2_outputs(1263)) xor (layer2_outputs(5817)));
    outputs(1510) <= layer2_outputs(9841);
    outputs(1511) <= not(layer2_outputs(7623));
    outputs(1512) <= layer2_outputs(10190);
    outputs(1513) <= not(layer2_outputs(8646));
    outputs(1514) <= (layer2_outputs(2823)) and not (layer2_outputs(1180));
    outputs(1515) <= (layer2_outputs(2503)) xor (layer2_outputs(2633));
    outputs(1516) <= not(layer2_outputs(5140));
    outputs(1517) <= not((layer2_outputs(6289)) xor (layer2_outputs(7072)));
    outputs(1518) <= layer2_outputs(550);
    outputs(1519) <= layer2_outputs(400);
    outputs(1520) <= (layer2_outputs(9431)) and not (layer2_outputs(3008));
    outputs(1521) <= (layer2_outputs(2989)) xor (layer2_outputs(9603));
    outputs(1522) <= not((layer2_outputs(3879)) xor (layer2_outputs(4619)));
    outputs(1523) <= layer2_outputs(10221);
    outputs(1524) <= (layer2_outputs(4699)) and (layer2_outputs(7355));
    outputs(1525) <= not(layer2_outputs(5065));
    outputs(1526) <= not((layer2_outputs(2412)) xor (layer2_outputs(4930)));
    outputs(1527) <= not((layer2_outputs(1621)) or (layer2_outputs(2935)));
    outputs(1528) <= layer2_outputs(6212);
    outputs(1529) <= not(layer2_outputs(1384));
    outputs(1530) <= not((layer2_outputs(2397)) xor (layer2_outputs(304)));
    outputs(1531) <= layer2_outputs(499);
    outputs(1532) <= (layer2_outputs(7899)) xor (layer2_outputs(445));
    outputs(1533) <= not((layer2_outputs(6171)) xor (layer2_outputs(3074)));
    outputs(1534) <= not((layer2_outputs(3306)) or (layer2_outputs(6869)));
    outputs(1535) <= layer2_outputs(4723);
    outputs(1536) <= (layer2_outputs(153)) and (layer2_outputs(3925));
    outputs(1537) <= not((layer2_outputs(2161)) or (layer2_outputs(8936)));
    outputs(1538) <= (layer2_outputs(7943)) and (layer2_outputs(4675));
    outputs(1539) <= not((layer2_outputs(7849)) xor (layer2_outputs(2107)));
    outputs(1540) <= (layer2_outputs(3278)) xor (layer2_outputs(9313));
    outputs(1541) <= (layer2_outputs(9112)) or (layer2_outputs(2167));
    outputs(1542) <= not((layer2_outputs(1474)) xor (layer2_outputs(6074)));
    outputs(1543) <= (layer2_outputs(8410)) xor (layer2_outputs(6202));
    outputs(1544) <= (layer2_outputs(7255)) xor (layer2_outputs(8455));
    outputs(1545) <= not(layer2_outputs(3594));
    outputs(1546) <= not((layer2_outputs(4676)) xor (layer2_outputs(9902)));
    outputs(1547) <= not((layer2_outputs(6854)) xor (layer2_outputs(7644)));
    outputs(1548) <= layer2_outputs(631);
    outputs(1549) <= (layer2_outputs(6751)) and not (layer2_outputs(2741));
    outputs(1550) <= layer2_outputs(1591);
    outputs(1551) <= (layer2_outputs(3834)) and (layer2_outputs(10094));
    outputs(1552) <= not(layer2_outputs(3448));
    outputs(1553) <= layer2_outputs(3858);
    outputs(1554) <= not(layer2_outputs(10079));
    outputs(1555) <= (layer2_outputs(8190)) and (layer2_outputs(996));
    outputs(1556) <= not((layer2_outputs(3540)) xor (layer2_outputs(3963)));
    outputs(1557) <= not((layer2_outputs(2564)) xor (layer2_outputs(914)));
    outputs(1558) <= layer2_outputs(7242);
    outputs(1559) <= not(layer2_outputs(6384)) or (layer2_outputs(4557));
    outputs(1560) <= not(layer2_outputs(8268));
    outputs(1561) <= not((layer2_outputs(5547)) xor (layer2_outputs(7836)));
    outputs(1562) <= not((layer2_outputs(5466)) xor (layer2_outputs(5646)));
    outputs(1563) <= (layer2_outputs(7672)) and (layer2_outputs(7889));
    outputs(1564) <= layer2_outputs(8538);
    outputs(1565) <= not((layer2_outputs(4001)) or (layer2_outputs(1935)));
    outputs(1566) <= (layer2_outputs(6363)) xor (layer2_outputs(823));
    outputs(1567) <= not((layer2_outputs(7736)) or (layer2_outputs(7)));
    outputs(1568) <= not((layer2_outputs(5815)) or (layer2_outputs(325)));
    outputs(1569) <= layer2_outputs(10117);
    outputs(1570) <= (layer2_outputs(1980)) xor (layer2_outputs(7739));
    outputs(1571) <= layer2_outputs(1053);
    outputs(1572) <= not((layer2_outputs(8882)) xor (layer2_outputs(10217)));
    outputs(1573) <= layer2_outputs(10086);
    outputs(1574) <= not(layer2_outputs(4470));
    outputs(1575) <= layer2_outputs(5239);
    outputs(1576) <= not(layer2_outputs(9498));
    outputs(1577) <= not(layer2_outputs(9157));
    outputs(1578) <= layer2_outputs(7074);
    outputs(1579) <= layer2_outputs(732);
    outputs(1580) <= not(layer2_outputs(5634));
    outputs(1581) <= (layer2_outputs(6396)) and not (layer2_outputs(3032));
    outputs(1582) <= not((layer2_outputs(9682)) or (layer2_outputs(1198)));
    outputs(1583) <= (layer2_outputs(6193)) xor (layer2_outputs(4497));
    outputs(1584) <= not((layer2_outputs(6722)) xor (layer2_outputs(6794)));
    outputs(1585) <= not(layer2_outputs(6501));
    outputs(1586) <= layer2_outputs(6158);
    outputs(1587) <= layer2_outputs(4861);
    outputs(1588) <= not(layer2_outputs(9946)) or (layer2_outputs(5586));
    outputs(1589) <= not(layer2_outputs(4649));
    outputs(1590) <= not((layer2_outputs(296)) or (layer2_outputs(6892)));
    outputs(1591) <= (layer2_outputs(7462)) and not (layer2_outputs(1228));
    outputs(1592) <= (layer2_outputs(6586)) xor (layer2_outputs(10229));
    outputs(1593) <= not(layer2_outputs(6978));
    outputs(1594) <= (layer2_outputs(3903)) or (layer2_outputs(6602));
    outputs(1595) <= not(layer2_outputs(5124));
    outputs(1596) <= (layer2_outputs(4017)) and not (layer2_outputs(7952));
    outputs(1597) <= (layer2_outputs(4474)) xor (layer2_outputs(688));
    outputs(1598) <= (layer2_outputs(2484)) xor (layer2_outputs(5001));
    outputs(1599) <= (layer2_outputs(6667)) xor (layer2_outputs(9589));
    outputs(1600) <= layer2_outputs(3821);
    outputs(1601) <= not((layer2_outputs(7194)) xor (layer2_outputs(8262)));
    outputs(1602) <= not((layer2_outputs(3455)) or (layer2_outputs(8388)));
    outputs(1603) <= not((layer2_outputs(2197)) xor (layer2_outputs(3931)));
    outputs(1604) <= layer2_outputs(7776);
    outputs(1605) <= not(layer2_outputs(1431));
    outputs(1606) <= not((layer2_outputs(1516)) and (layer2_outputs(5498)));
    outputs(1607) <= not((layer2_outputs(8440)) xor (layer2_outputs(3369)));
    outputs(1608) <= layer2_outputs(3792);
    outputs(1609) <= (layer2_outputs(4890)) and not (layer2_outputs(2844));
    outputs(1610) <= (layer2_outputs(3598)) and not (layer2_outputs(670));
    outputs(1611) <= not(layer2_outputs(5374));
    outputs(1612) <= layer2_outputs(5340);
    outputs(1613) <= not((layer2_outputs(435)) xor (layer2_outputs(7358)));
    outputs(1614) <= layer2_outputs(3705);
    outputs(1615) <= not(layer2_outputs(3309));
    outputs(1616) <= (layer2_outputs(453)) xor (layer2_outputs(6956));
    outputs(1617) <= not(layer2_outputs(1185));
    outputs(1618) <= not((layer2_outputs(8322)) or (layer2_outputs(3454)));
    outputs(1619) <= not(layer2_outputs(5020));
    outputs(1620) <= (layer2_outputs(1445)) and not (layer2_outputs(6653));
    outputs(1621) <= layer2_outputs(9983);
    outputs(1622) <= not((layer2_outputs(3434)) xor (layer2_outputs(9743)));
    outputs(1623) <= (layer2_outputs(356)) xor (layer2_outputs(3204));
    outputs(1624) <= layer2_outputs(3385);
    outputs(1625) <= not(layer2_outputs(5828));
    outputs(1626) <= (layer2_outputs(5640)) and not (layer2_outputs(7507));
    outputs(1627) <= not((layer2_outputs(5021)) xor (layer2_outputs(2902)));
    outputs(1628) <= not((layer2_outputs(3917)) xor (layer2_outputs(1108)));
    outputs(1629) <= (layer2_outputs(3204)) and (layer2_outputs(518));
    outputs(1630) <= not(layer2_outputs(7713));
    outputs(1631) <= layer2_outputs(7556);
    outputs(1632) <= not((layer2_outputs(3740)) or (layer2_outputs(1103)));
    outputs(1633) <= not((layer2_outputs(7997)) xor (layer2_outputs(3610)));
    outputs(1634) <= layer2_outputs(9529);
    outputs(1635) <= (layer2_outputs(6241)) and not (layer2_outputs(5892));
    outputs(1636) <= not(layer2_outputs(7198));
    outputs(1637) <= layer2_outputs(2558);
    outputs(1638) <= (layer2_outputs(2979)) xor (layer2_outputs(6449));
    outputs(1639) <= (layer2_outputs(5619)) and not (layer2_outputs(3231));
    outputs(1640) <= (layer2_outputs(5799)) and not (layer2_outputs(7731));
    outputs(1641) <= (layer2_outputs(8726)) xor (layer2_outputs(3667));
    outputs(1642) <= not(layer2_outputs(4223)) or (layer2_outputs(8520));
    outputs(1643) <= not((layer2_outputs(8093)) xor (layer2_outputs(8085)));
    outputs(1644) <= layer2_outputs(2960);
    outputs(1645) <= (layer2_outputs(4766)) and (layer2_outputs(879));
    outputs(1646) <= not((layer2_outputs(4385)) xor (layer2_outputs(6563)));
    outputs(1647) <= not(layer2_outputs(1464));
    outputs(1648) <= not((layer2_outputs(1445)) xor (layer2_outputs(9306)));
    outputs(1649) <= not(layer2_outputs(9262));
    outputs(1650) <= (layer2_outputs(7655)) xor (layer2_outputs(9729));
    outputs(1651) <= (layer2_outputs(9248)) xor (layer2_outputs(4704));
    outputs(1652) <= (layer2_outputs(8362)) and not (layer2_outputs(3046));
    outputs(1653) <= layer2_outputs(5477);
    outputs(1654) <= (layer2_outputs(759)) xor (layer2_outputs(6861));
    outputs(1655) <= (layer2_outputs(10227)) and not (layer2_outputs(5071));
    outputs(1656) <= not((layer2_outputs(8258)) or (layer2_outputs(1278)));
    outputs(1657) <= layer2_outputs(6317);
    outputs(1658) <= layer2_outputs(3755);
    outputs(1659) <= not((layer2_outputs(7188)) xor (layer2_outputs(413)));
    outputs(1660) <= not(layer2_outputs(5351));
    outputs(1661) <= not(layer2_outputs(289));
    outputs(1662) <= (layer2_outputs(3724)) and not (layer2_outputs(3198));
    outputs(1663) <= layer2_outputs(3498);
    outputs(1664) <= (layer2_outputs(7989)) and (layer2_outputs(440));
    outputs(1665) <= not(layer2_outputs(9930));
    outputs(1666) <= layer2_outputs(5133);
    outputs(1667) <= not((layer2_outputs(5592)) xor (layer2_outputs(643)));
    outputs(1668) <= layer2_outputs(10060);
    outputs(1669) <= layer2_outputs(1592);
    outputs(1670) <= not((layer2_outputs(4549)) xor (layer2_outputs(6455)));
    outputs(1671) <= (layer2_outputs(365)) and not (layer2_outputs(2143));
    outputs(1672) <= layer2_outputs(4722);
    outputs(1673) <= layer2_outputs(710);
    outputs(1674) <= not((layer2_outputs(7950)) xor (layer2_outputs(4690)));
    outputs(1675) <= layer2_outputs(7008);
    outputs(1676) <= not(layer2_outputs(4353));
    outputs(1677) <= not(layer2_outputs(5380));
    outputs(1678) <= layer2_outputs(518);
    outputs(1679) <= not((layer2_outputs(1748)) xor (layer2_outputs(446)));
    outputs(1680) <= not((layer2_outputs(7475)) and (layer2_outputs(7848)));
    outputs(1681) <= (layer2_outputs(5307)) and (layer2_outputs(3440));
    outputs(1682) <= (layer2_outputs(5485)) xor (layer2_outputs(4651));
    outputs(1683) <= (layer2_outputs(7108)) and not (layer2_outputs(4898));
    outputs(1684) <= (layer2_outputs(800)) xor (layer2_outputs(8707));
    outputs(1685) <= not(layer2_outputs(2123));
    outputs(1686) <= (layer2_outputs(9003)) and (layer2_outputs(7944));
    outputs(1687) <= not(layer2_outputs(10137));
    outputs(1688) <= (layer2_outputs(8083)) xor (layer2_outputs(2205));
    outputs(1689) <= layer2_outputs(5627);
    outputs(1690) <= (layer2_outputs(8180)) xor (layer2_outputs(6181));
    outputs(1691) <= not((layer2_outputs(2347)) xor (layer2_outputs(6893)));
    outputs(1692) <= not(layer2_outputs(1123));
    outputs(1693) <= (layer2_outputs(8302)) xor (layer2_outputs(5795));
    outputs(1694) <= layer2_outputs(8153);
    outputs(1695) <= layer2_outputs(8401);
    outputs(1696) <= layer2_outputs(310);
    outputs(1697) <= not(layer2_outputs(3487)) or (layer2_outputs(6381));
    outputs(1698) <= not((layer2_outputs(3263)) or (layer2_outputs(5656)));
    outputs(1699) <= layer2_outputs(3929);
    outputs(1700) <= not((layer2_outputs(9374)) xor (layer2_outputs(5559)));
    outputs(1701) <= (layer2_outputs(1042)) and (layer2_outputs(5572));
    outputs(1702) <= not((layer2_outputs(4989)) xor (layer2_outputs(1060)));
    outputs(1703) <= not((layer2_outputs(7901)) xor (layer2_outputs(4449)));
    outputs(1704) <= (layer2_outputs(2168)) and (layer2_outputs(10));
    outputs(1705) <= not((layer2_outputs(9620)) xor (layer2_outputs(5650)));
    outputs(1706) <= layer2_outputs(8032);
    outputs(1707) <= layer2_outputs(9993);
    outputs(1708) <= not((layer2_outputs(4733)) or (layer2_outputs(66)));
    outputs(1709) <= (layer2_outputs(4193)) and not (layer2_outputs(6964));
    outputs(1710) <= (layer2_outputs(7291)) xor (layer2_outputs(1834));
    outputs(1711) <= (layer2_outputs(479)) and not (layer2_outputs(7373));
    outputs(1712) <= not((layer2_outputs(752)) xor (layer2_outputs(1296)));
    outputs(1713) <= (layer2_outputs(10212)) xor (layer2_outputs(628));
    outputs(1714) <= not(layer2_outputs(6898));
    outputs(1715) <= not(layer2_outputs(2680));
    outputs(1716) <= layer2_outputs(1092);
    outputs(1717) <= not(layer2_outputs(4114)) or (layer2_outputs(6558));
    outputs(1718) <= layer2_outputs(9865);
    outputs(1719) <= layer2_outputs(5989);
    outputs(1720) <= not((layer2_outputs(1640)) or (layer2_outputs(9166)));
    outputs(1721) <= layer2_outputs(3849);
    outputs(1722) <= (layer2_outputs(2298)) xor (layer2_outputs(9163));
    outputs(1723) <= not(layer2_outputs(1291));
    outputs(1724) <= (layer2_outputs(7893)) and not (layer2_outputs(7168));
    outputs(1725) <= not(layer2_outputs(9033));
    outputs(1726) <= not((layer2_outputs(6172)) xor (layer2_outputs(1484)));
    outputs(1727) <= layer2_outputs(6134);
    outputs(1728) <= layer2_outputs(923);
    outputs(1729) <= (layer2_outputs(357)) xor (layer2_outputs(3891));
    outputs(1730) <= not((layer2_outputs(6488)) xor (layer2_outputs(7204)));
    outputs(1731) <= (layer2_outputs(7298)) xor (layer2_outputs(2807));
    outputs(1732) <= (layer2_outputs(2162)) xor (layer2_outputs(4599));
    outputs(1733) <= layer2_outputs(8000);
    outputs(1734) <= not((layer2_outputs(4440)) xor (layer2_outputs(6655)));
    outputs(1735) <= not(layer2_outputs(5285));
    outputs(1736) <= (layer2_outputs(3030)) and (layer2_outputs(8698));
    outputs(1737) <= not((layer2_outputs(3216)) xor (layer2_outputs(6504)));
    outputs(1738) <= not(layer2_outputs(1226));
    outputs(1739) <= not(layer2_outputs(2507)) or (layer2_outputs(8481));
    outputs(1740) <= not(layer2_outputs(5444));
    outputs(1741) <= layer2_outputs(4220);
    outputs(1742) <= not((layer2_outputs(3309)) and (layer2_outputs(8335)));
    outputs(1743) <= not((layer2_outputs(2478)) or (layer2_outputs(4572)));
    outputs(1744) <= not(layer2_outputs(4775));
    outputs(1745) <= layer2_outputs(5658);
    outputs(1746) <= layer2_outputs(9212);
    outputs(1747) <= layer2_outputs(1982);
    outputs(1748) <= (layer2_outputs(9529)) or (layer2_outputs(9072));
    outputs(1749) <= not(layer2_outputs(4046));
    outputs(1750) <= (layer2_outputs(2510)) and not (layer2_outputs(3478));
    outputs(1751) <= layer2_outputs(4044);
    outputs(1752) <= not(layer2_outputs(1876));
    outputs(1753) <= not((layer2_outputs(2405)) and (layer2_outputs(3468)));
    outputs(1754) <= not((layer2_outputs(469)) and (layer2_outputs(5773)));
    outputs(1755) <= not(layer2_outputs(4043));
    outputs(1756) <= layer2_outputs(1897);
    outputs(1757) <= not(layer2_outputs(9116));
    outputs(1758) <= not(layer2_outputs(4480));
    outputs(1759) <= not((layer2_outputs(5868)) xor (layer2_outputs(2383)));
    outputs(1760) <= (layer2_outputs(3176)) xor (layer2_outputs(1294));
    outputs(1761) <= (layer2_outputs(419)) xor (layer2_outputs(1231));
    outputs(1762) <= not(layer2_outputs(3288));
    outputs(1763) <= (layer2_outputs(3975)) and not (layer2_outputs(5493));
    outputs(1764) <= (layer2_outputs(8954)) and not (layer2_outputs(6636));
    outputs(1765) <= not((layer2_outputs(7547)) xor (layer2_outputs(6326)));
    outputs(1766) <= not(layer2_outputs(6848));
    outputs(1767) <= not((layer2_outputs(7655)) xor (layer2_outputs(5286)));
    outputs(1768) <= not((layer2_outputs(302)) xor (layer2_outputs(7860)));
    outputs(1769) <= not((layer2_outputs(9081)) and (layer2_outputs(6870)));
    outputs(1770) <= layer2_outputs(2843);
    outputs(1771) <= not(layer2_outputs(3690));
    outputs(1772) <= (layer2_outputs(6854)) xor (layer2_outputs(7645));
    outputs(1773) <= (layer2_outputs(3556)) and (layer2_outputs(2963));
    outputs(1774) <= (layer2_outputs(4860)) xor (layer2_outputs(2783));
    outputs(1775) <= not((layer2_outputs(8885)) or (layer2_outputs(3599)));
    outputs(1776) <= (layer2_outputs(9613)) and not (layer2_outputs(10138));
    outputs(1777) <= (layer2_outputs(4148)) and not (layer2_outputs(5793));
    outputs(1778) <= not((layer2_outputs(6367)) or (layer2_outputs(6067)));
    outputs(1779) <= (layer2_outputs(9875)) and not (layer2_outputs(2296));
    outputs(1780) <= not(layer2_outputs(1436));
    outputs(1781) <= (layer2_outputs(1062)) xor (layer2_outputs(1598));
    outputs(1782) <= (layer2_outputs(8672)) xor (layer2_outputs(7402));
    outputs(1783) <= not(layer2_outputs(6863));
    outputs(1784) <= layer2_outputs(9089);
    outputs(1785) <= (layer2_outputs(7770)) and not (layer2_outputs(2346));
    outputs(1786) <= (layer2_outputs(4231)) and not (layer2_outputs(5471));
    outputs(1787) <= (layer2_outputs(3897)) and not (layer2_outputs(8431));
    outputs(1788) <= layer2_outputs(9168);
    outputs(1789) <= not((layer2_outputs(777)) xor (layer2_outputs(3871)));
    outputs(1790) <= (layer2_outputs(8594)) and not (layer2_outputs(6678));
    outputs(1791) <= layer2_outputs(8434);
    outputs(1792) <= not(layer2_outputs(846));
    outputs(1793) <= not(layer2_outputs(6975));
    outputs(1794) <= (layer2_outputs(6980)) and not (layer2_outputs(972));
    outputs(1795) <= not(layer2_outputs(6979));
    outputs(1796) <= layer2_outputs(3460);
    outputs(1797) <= layer2_outputs(8237);
    outputs(1798) <= not(layer2_outputs(9424));
    outputs(1799) <= layer2_outputs(6275);
    outputs(1800) <= (layer2_outputs(6608)) xor (layer2_outputs(6904));
    outputs(1801) <= (layer2_outputs(2232)) and not (layer2_outputs(1704));
    outputs(1802) <= (layer2_outputs(1170)) and not (layer2_outputs(481));
    outputs(1803) <= not(layer2_outputs(4984));
    outputs(1804) <= not((layer2_outputs(1908)) or (layer2_outputs(6081)));
    outputs(1805) <= not(layer2_outputs(9207));
    outputs(1806) <= not((layer2_outputs(7224)) or (layer2_outputs(8039)));
    outputs(1807) <= not((layer2_outputs(4833)) xor (layer2_outputs(5161)));
    outputs(1808) <= not((layer2_outputs(260)) or (layer2_outputs(6352)));
    outputs(1809) <= layer2_outputs(8531);
    outputs(1810) <= not(layer2_outputs(2918));
    outputs(1811) <= layer2_outputs(7462);
    outputs(1812) <= layer2_outputs(5047);
    outputs(1813) <= not(layer2_outputs(5403));
    outputs(1814) <= not(layer2_outputs(7139));
    outputs(1815) <= (layer2_outputs(6730)) and not (layer2_outputs(3547));
    outputs(1816) <= (layer2_outputs(2286)) and not (layer2_outputs(5389));
    outputs(1817) <= layer2_outputs(7708);
    outputs(1818) <= not(layer2_outputs(5363)) or (layer2_outputs(3966));
    outputs(1819) <= (layer2_outputs(6140)) and not (layer2_outputs(9405));
    outputs(1820) <= layer2_outputs(8701);
    outputs(1821) <= not((layer2_outputs(7347)) or (layer2_outputs(2802)));
    outputs(1822) <= layer2_outputs(9181);
    outputs(1823) <= (layer2_outputs(7465)) and (layer2_outputs(8992));
    outputs(1824) <= not((layer2_outputs(4762)) xor (layer2_outputs(7292)));
    outputs(1825) <= (layer2_outputs(3234)) xor (layer2_outputs(330));
    outputs(1826) <= layer2_outputs(7166);
    outputs(1827) <= not((layer2_outputs(2985)) or (layer2_outputs(6522)));
    outputs(1828) <= (layer2_outputs(8958)) xor (layer2_outputs(5874));
    outputs(1829) <= not((layer2_outputs(4907)) or (layer2_outputs(1131)));
    outputs(1830) <= not(layer2_outputs(5064));
    outputs(1831) <= not(layer2_outputs(7949));
    outputs(1832) <= layer2_outputs(9565);
    outputs(1833) <= not(layer2_outputs(4199));
    outputs(1834) <= '0';
    outputs(1835) <= (layer2_outputs(8270)) and not (layer2_outputs(5083));
    outputs(1836) <= (layer2_outputs(8657)) xor (layer2_outputs(4014));
    outputs(1837) <= not((layer2_outputs(1253)) xor (layer2_outputs(363)));
    outputs(1838) <= not(layer2_outputs(5331)) or (layer2_outputs(4039));
    outputs(1839) <= (layer2_outputs(9504)) and (layer2_outputs(641));
    outputs(1840) <= layer2_outputs(7974);
    outputs(1841) <= not((layer2_outputs(5537)) or (layer2_outputs(266)));
    outputs(1842) <= not(layer2_outputs(7104));
    outputs(1843) <= layer2_outputs(5971);
    outputs(1844) <= not(layer2_outputs(9674));
    outputs(1845) <= not((layer2_outputs(8737)) and (layer2_outputs(7070)));
    outputs(1846) <= layer2_outputs(3459);
    outputs(1847) <= (layer2_outputs(141)) xor (layer2_outputs(769));
    outputs(1848) <= (layer2_outputs(7309)) and (layer2_outputs(5143));
    outputs(1849) <= (layer2_outputs(673)) and not (layer2_outputs(4604));
    outputs(1850) <= not(layer2_outputs(4466));
    outputs(1851) <= not((layer2_outputs(5420)) xor (layer2_outputs(8386)));
    outputs(1852) <= not((layer2_outputs(7878)) or (layer2_outputs(8428)));
    outputs(1853) <= not((layer2_outputs(329)) or (layer2_outputs(4649)));
    outputs(1854) <= not((layer2_outputs(761)) xor (layer2_outputs(1213)));
    outputs(1855) <= (layer2_outputs(7687)) xor (layer2_outputs(5255));
    outputs(1856) <= (layer2_outputs(5961)) and (layer2_outputs(6036));
    outputs(1857) <= layer2_outputs(7922);
    outputs(1858) <= not(layer2_outputs(6930));
    outputs(1859) <= (layer2_outputs(8697)) and not (layer2_outputs(9847));
    outputs(1860) <= (layer2_outputs(3542)) xor (layer2_outputs(7500));
    outputs(1861) <= not((layer2_outputs(6699)) or (layer2_outputs(84)));
    outputs(1862) <= (layer2_outputs(6487)) xor (layer2_outputs(1676));
    outputs(1863) <= not(layer2_outputs(9321));
    outputs(1864) <= layer2_outputs(6663);
    outputs(1865) <= (layer2_outputs(3631)) and not (layer2_outputs(530));
    outputs(1866) <= not((layer2_outputs(2794)) xor (layer2_outputs(9173)));
    outputs(1867) <= not((layer2_outputs(9882)) xor (layer2_outputs(2118)));
    outputs(1868) <= (layer2_outputs(4573)) xor (layer2_outputs(5932));
    outputs(1869) <= (layer2_outputs(1003)) xor (layer2_outputs(2224));
    outputs(1870) <= layer2_outputs(67);
    outputs(1871) <= (layer2_outputs(7304)) and (layer2_outputs(1288));
    outputs(1872) <= layer2_outputs(4507);
    outputs(1873) <= not((layer2_outputs(5337)) xor (layer2_outputs(9414)));
    outputs(1874) <= not(layer2_outputs(3310));
    outputs(1875) <= (layer2_outputs(5891)) and not (layer2_outputs(2764));
    outputs(1876) <= (layer2_outputs(9369)) and (layer2_outputs(6354));
    outputs(1877) <= not(layer2_outputs(3117));
    outputs(1878) <= (layer2_outputs(8353)) xor (layer2_outputs(4257));
    outputs(1879) <= (layer2_outputs(6329)) and (layer2_outputs(8827));
    outputs(1880) <= (layer2_outputs(33)) and not (layer2_outputs(8503));
    outputs(1881) <= not(layer2_outputs(1789));
    outputs(1882) <= not(layer2_outputs(2899));
    outputs(1883) <= not(layer2_outputs(5381));
    outputs(1884) <= (layer2_outputs(9557)) xor (layer2_outputs(4730));
    outputs(1885) <= not(layer2_outputs(823)) or (layer2_outputs(4797));
    outputs(1886) <= not(layer2_outputs(9146));
    outputs(1887) <= (layer2_outputs(6832)) and not (layer2_outputs(5093));
    outputs(1888) <= layer2_outputs(3226);
    outputs(1889) <= not(layer2_outputs(3513));
    outputs(1890) <= not((layer2_outputs(4647)) xor (layer2_outputs(3101)));
    outputs(1891) <= (layer2_outputs(9899)) and (layer2_outputs(232));
    outputs(1892) <= not(layer2_outputs(6343));
    outputs(1893) <= layer2_outputs(3884);
    outputs(1894) <= layer2_outputs(9765);
    outputs(1895) <= (layer2_outputs(7865)) xor (layer2_outputs(2654));
    outputs(1896) <= (layer2_outputs(2394)) and not (layer2_outputs(10139));
    outputs(1897) <= not(layer2_outputs(9956));
    outputs(1898) <= (layer2_outputs(4987)) and (layer2_outputs(2871));
    outputs(1899) <= (layer2_outputs(4735)) and (layer2_outputs(7489));
    outputs(1900) <= not((layer2_outputs(7025)) xor (layer2_outputs(7808)));
    outputs(1901) <= not((layer2_outputs(3095)) xor (layer2_outputs(6908)));
    outputs(1902) <= (layer2_outputs(5798)) and not (layer2_outputs(598));
    outputs(1903) <= (layer2_outputs(10114)) xor (layer2_outputs(74));
    outputs(1904) <= not((layer2_outputs(4904)) or (layer2_outputs(793)));
    outputs(1905) <= not((layer2_outputs(617)) xor (layer2_outputs(5473)));
    outputs(1906) <= (layer2_outputs(3301)) and not (layer2_outputs(3655));
    outputs(1907) <= not((layer2_outputs(980)) xor (layer2_outputs(4924)));
    outputs(1908) <= not((layer2_outputs(3816)) or (layer2_outputs(4263)));
    outputs(1909) <= not(layer2_outputs(3201));
    outputs(1910) <= (layer2_outputs(2690)) and (layer2_outputs(698));
    outputs(1911) <= layer2_outputs(8359);
    outputs(1912) <= not((layer2_outputs(5433)) xor (layer2_outputs(9218)));
    outputs(1913) <= (layer2_outputs(325)) xor (layer2_outputs(8998));
    outputs(1914) <= (layer2_outputs(3189)) and (layer2_outputs(1840));
    outputs(1915) <= (layer2_outputs(4002)) and not (layer2_outputs(2940));
    outputs(1916) <= (layer2_outputs(7972)) and not (layer2_outputs(9770));
    outputs(1917) <= (layer2_outputs(4666)) and not (layer2_outputs(9888));
    outputs(1918) <= (layer2_outputs(6651)) xor (layer2_outputs(2142));
    outputs(1919) <= not(layer2_outputs(4150));
    outputs(1920) <= layer2_outputs(5232);
    outputs(1921) <= not((layer2_outputs(9789)) xor (layer2_outputs(4577)));
    outputs(1922) <= not(layer2_outputs(7018));
    outputs(1923) <= not(layer2_outputs(7935));
    outputs(1924) <= not((layer2_outputs(2282)) xor (layer2_outputs(8290)));
    outputs(1925) <= not(layer2_outputs(4732));
    outputs(1926) <= (layer2_outputs(7491)) xor (layer2_outputs(3062));
    outputs(1927) <= not(layer2_outputs(9619));
    outputs(1928) <= layer2_outputs(3160);
    outputs(1929) <= layer2_outputs(4401);
    outputs(1930) <= not(layer2_outputs(1912));
    outputs(1931) <= not(layer2_outputs(5858));
    outputs(1932) <= (layer2_outputs(2821)) xor (layer2_outputs(1168));
    outputs(1933) <= (layer2_outputs(3774)) xor (layer2_outputs(3940));
    outputs(1934) <= '0';
    outputs(1935) <= not(layer2_outputs(5224));
    outputs(1936) <= not((layer2_outputs(4606)) xor (layer2_outputs(9631)));
    outputs(1937) <= not((layer2_outputs(6963)) xor (layer2_outputs(5106)));
    outputs(1938) <= layer2_outputs(4190);
    outputs(1939) <= (layer2_outputs(2999)) and not (layer2_outputs(4772));
    outputs(1940) <= (layer2_outputs(6329)) and not (layer2_outputs(9997));
    outputs(1941) <= layer2_outputs(2849);
    outputs(1942) <= (layer2_outputs(8632)) and not (layer2_outputs(991));
    outputs(1943) <= layer2_outputs(9611);
    outputs(1944) <= not(layer2_outputs(9805));
    outputs(1945) <= not((layer2_outputs(5556)) or (layer2_outputs(4462)));
    outputs(1946) <= not(layer2_outputs(8646));
    outputs(1947) <= not((layer2_outputs(6612)) or (layer2_outputs(410)));
    outputs(1948) <= not((layer2_outputs(4899)) xor (layer2_outputs(3823)));
    outputs(1949) <= not((layer2_outputs(3077)) xor (layer2_outputs(8630)));
    outputs(1950) <= not(layer2_outputs(1669));
    outputs(1951) <= (layer2_outputs(7206)) and not (layer2_outputs(9397));
    outputs(1952) <= not(layer2_outputs(492));
    outputs(1953) <= not(layer2_outputs(4457));
    outputs(1954) <= not(layer2_outputs(1887));
    outputs(1955) <= not(layer2_outputs(2459));
    outputs(1956) <= not(layer2_outputs(9289));
    outputs(1957) <= not((layer2_outputs(1889)) xor (layer2_outputs(4716)));
    outputs(1958) <= not((layer2_outputs(4502)) or (layer2_outputs(1376)));
    outputs(1959) <= (layer2_outputs(1284)) and (layer2_outputs(9648));
    outputs(1960) <= not(layer2_outputs(7055));
    outputs(1961) <= not((layer2_outputs(1626)) xor (layer2_outputs(557)));
    outputs(1962) <= not((layer2_outputs(3742)) xor (layer2_outputs(7199)));
    outputs(1963) <= (layer2_outputs(8316)) and not (layer2_outputs(195));
    outputs(1964) <= (layer2_outputs(2144)) and not (layer2_outputs(7316));
    outputs(1965) <= layer2_outputs(2208);
    outputs(1966) <= not(layer2_outputs(6286));
    outputs(1967) <= not(layer2_outputs(7335));
    outputs(1968) <= (layer2_outputs(474)) and not (layer2_outputs(943));
    outputs(1969) <= layer2_outputs(9843);
    outputs(1970) <= not(layer2_outputs(1369));
    outputs(1971) <= '0';
    outputs(1972) <= layer2_outputs(5711);
    outputs(1973) <= not(layer2_outputs(4098));
    outputs(1974) <= layer2_outputs(7484);
    outputs(1975) <= layer2_outputs(4476);
    outputs(1976) <= not((layer2_outputs(4054)) xor (layer2_outputs(8172)));
    outputs(1977) <= not(layer2_outputs(1539));
    outputs(1978) <= not(layer2_outputs(2227));
    outputs(1979) <= (layer2_outputs(1850)) and not (layer2_outputs(1427));
    outputs(1980) <= (layer2_outputs(5223)) and not (layer2_outputs(3646));
    outputs(1981) <= not(layer2_outputs(177));
    outputs(1982) <= layer2_outputs(167);
    outputs(1983) <= (layer2_outputs(7544)) xor (layer2_outputs(5754));
    outputs(1984) <= not((layer2_outputs(4593)) xor (layer2_outputs(8655)));
    outputs(1985) <= layer2_outputs(6053);
    outputs(1986) <= not(layer2_outputs(2573));
    outputs(1987) <= layer2_outputs(3618);
    outputs(1988) <= (layer2_outputs(7324)) xor (layer2_outputs(7411));
    outputs(1989) <= not(layer2_outputs(8647));
    outputs(1990) <= (layer2_outputs(2922)) and not (layer2_outputs(4032));
    outputs(1991) <= layer2_outputs(2811);
    outputs(1992) <= (layer2_outputs(4546)) and (layer2_outputs(3187));
    outputs(1993) <= not(layer2_outputs(1123));
    outputs(1994) <= not(layer2_outputs(8535));
    outputs(1995) <= layer2_outputs(2074);
    outputs(1996) <= not((layer2_outputs(8920)) xor (layer2_outputs(858)));
    outputs(1997) <= not(layer2_outputs(1690));
    outputs(1998) <= '0';
    outputs(1999) <= not(layer2_outputs(7103));
    outputs(2000) <= not((layer2_outputs(7144)) xor (layer2_outputs(2883)));
    outputs(2001) <= (layer2_outputs(10197)) xor (layer2_outputs(4645));
    outputs(2002) <= layer2_outputs(5030);
    outputs(2003) <= not((layer2_outputs(1407)) xor (layer2_outputs(394)));
    outputs(2004) <= layer2_outputs(4908);
    outputs(2005) <= not((layer2_outputs(5147)) or (layer2_outputs(9515)));
    outputs(2006) <= (layer2_outputs(9023)) and (layer2_outputs(5343));
    outputs(2007) <= not(layer2_outputs(6520));
    outputs(2008) <= not((layer2_outputs(7582)) xor (layer2_outputs(3713)));
    outputs(2009) <= layer2_outputs(3506);
    outputs(2010) <= (layer2_outputs(1352)) and (layer2_outputs(2761));
    outputs(2011) <= not((layer2_outputs(3516)) xor (layer2_outputs(8647)));
    outputs(2012) <= not((layer2_outputs(8029)) xor (layer2_outputs(948)));
    outputs(2013) <= not(layer2_outputs(9193));
    outputs(2014) <= layer2_outputs(1158);
    outputs(2015) <= not((layer2_outputs(7819)) xor (layer2_outputs(8044)));
    outputs(2016) <= not(layer2_outputs(2717));
    outputs(2017) <= (layer2_outputs(6714)) and not (layer2_outputs(7754));
    outputs(2018) <= layer2_outputs(2626);
    outputs(2019) <= not((layer2_outputs(6226)) xor (layer2_outputs(7648)));
    outputs(2020) <= layer2_outputs(3264);
    outputs(2021) <= (layer2_outputs(6937)) and not (layer2_outputs(6998));
    outputs(2022) <= (layer2_outputs(6794)) xor (layer2_outputs(1739));
    outputs(2023) <= not((layer2_outputs(5875)) xor (layer2_outputs(4437)));
    outputs(2024) <= layer2_outputs(5376);
    outputs(2025) <= not(layer2_outputs(5497));
    outputs(2026) <= (layer2_outputs(5971)) and not (layer2_outputs(3070));
    outputs(2027) <= '0';
    outputs(2028) <= not((layer2_outputs(3530)) or (layer2_outputs(4586)));
    outputs(2029) <= not(layer2_outputs(2278));
    outputs(2030) <= layer2_outputs(7115);
    outputs(2031) <= layer2_outputs(10099);
    outputs(2032) <= (layer2_outputs(7756)) xor (layer2_outputs(6784));
    outputs(2033) <= not(layer2_outputs(5356));
    outputs(2034) <= not(layer2_outputs(6631));
    outputs(2035) <= (layer2_outputs(441)) and not (layer2_outputs(8663));
    outputs(2036) <= layer2_outputs(5000);
    outputs(2037) <= layer2_outputs(5171);
    outputs(2038) <= not(layer2_outputs(403));
    outputs(2039) <= (layer2_outputs(4544)) xor (layer2_outputs(8696));
    outputs(2040) <= not((layer2_outputs(9697)) xor (layer2_outputs(5522)));
    outputs(2041) <= not(layer2_outputs(41));
    outputs(2042) <= layer2_outputs(1710);
    outputs(2043) <= not(layer2_outputs(241));
    outputs(2044) <= not(layer2_outputs(6913));
    outputs(2045) <= not((layer2_outputs(7155)) xor (layer2_outputs(7663)));
    outputs(2046) <= (layer2_outputs(6754)) and (layer2_outputs(1435));
    outputs(2047) <= (layer2_outputs(8203)) xor (layer2_outputs(2949));
    outputs(2048) <= not((layer2_outputs(1702)) or (layer2_outputs(3652)));
    outputs(2049) <= not((layer2_outputs(9653)) and (layer2_outputs(5088)));
    outputs(2050) <= not(layer2_outputs(4284));
    outputs(2051) <= (layer2_outputs(2209)) and (layer2_outputs(707));
    outputs(2052) <= layer2_outputs(1751);
    outputs(2053) <= not(layer2_outputs(9808));
    outputs(2054) <= layer2_outputs(4230);
    outputs(2055) <= layer2_outputs(8533);
    outputs(2056) <= layer2_outputs(7791);
    outputs(2057) <= not((layer2_outputs(2354)) or (layer2_outputs(5012)));
    outputs(2058) <= layer2_outputs(9967);
    outputs(2059) <= (layer2_outputs(8880)) xor (layer2_outputs(2788));
    outputs(2060) <= not((layer2_outputs(10039)) and (layer2_outputs(9331)));
    outputs(2061) <= not(layer2_outputs(6922));
    outputs(2062) <= layer2_outputs(194);
    outputs(2063) <= not(layer2_outputs(6685));
    outputs(2064) <= not(layer2_outputs(5731)) or (layer2_outputs(844));
    outputs(2065) <= not((layer2_outputs(7961)) xor (layer2_outputs(1139)));
    outputs(2066) <= not(layer2_outputs(4253));
    outputs(2067) <= not(layer2_outputs(6339));
    outputs(2068) <= not(layer2_outputs(3413)) or (layer2_outputs(5780));
    outputs(2069) <= layer2_outputs(9476);
    outputs(2070) <= layer2_outputs(4958);
    outputs(2071) <= not(layer2_outputs(816)) or (layer2_outputs(2702));
    outputs(2072) <= not(layer2_outputs(3714));
    outputs(2073) <= layer2_outputs(788);
    outputs(2074) <= not(layer2_outputs(9665));
    outputs(2075) <= not((layer2_outputs(1450)) or (layer2_outputs(9743)));
    outputs(2076) <= layer2_outputs(61);
    outputs(2077) <= not(layer2_outputs(122));
    outputs(2078) <= (layer2_outputs(2740)) xor (layer2_outputs(924));
    outputs(2079) <= layer2_outputs(1922);
    outputs(2080) <= layer2_outputs(3171);
    outputs(2081) <= not((layer2_outputs(2055)) and (layer2_outputs(3669)));
    outputs(2082) <= layer2_outputs(5066);
    outputs(2083) <= layer2_outputs(6737);
    outputs(2084) <= not((layer2_outputs(8819)) or (layer2_outputs(4033)));
    outputs(2085) <= not(layer2_outputs(6641));
    outputs(2086) <= not((layer2_outputs(9240)) or (layer2_outputs(3410)));
    outputs(2087) <= not((layer2_outputs(2106)) xor (layer2_outputs(5378)));
    outputs(2088) <= layer2_outputs(10141);
    outputs(2089) <= not(layer2_outputs(5900));
    outputs(2090) <= (layer2_outputs(7771)) and not (layer2_outputs(10025));
    outputs(2091) <= not((layer2_outputs(4421)) and (layer2_outputs(3545)));
    outputs(2092) <= not(layer2_outputs(4108));
    outputs(2093) <= not((layer2_outputs(634)) xor (layer2_outputs(4327)));
    outputs(2094) <= layer2_outputs(9481);
    outputs(2095) <= layer2_outputs(2694);
    outputs(2096) <= not((layer2_outputs(6632)) xor (layer2_outputs(5620)));
    outputs(2097) <= not(layer2_outputs(6090)) or (layer2_outputs(4935));
    outputs(2098) <= layer2_outputs(6977);
    outputs(2099) <= (layer2_outputs(1262)) and not (layer2_outputs(2163));
    outputs(2100) <= (layer2_outputs(2411)) and not (layer2_outputs(7996));
    outputs(2101) <= not(layer2_outputs(5192));
    outputs(2102) <= (layer2_outputs(8202)) xor (layer2_outputs(859));
    outputs(2103) <= not(layer2_outputs(1232));
    outputs(2104) <= layer2_outputs(4436);
    outputs(2105) <= layer2_outputs(5207);
    outputs(2106) <= layer2_outputs(3201);
    outputs(2107) <= not(layer2_outputs(3743));
    outputs(2108) <= layer2_outputs(2254);
    outputs(2109) <= (layer2_outputs(4004)) and not (layer2_outputs(6503));
    outputs(2110) <= layer2_outputs(1361);
    outputs(2111) <= layer2_outputs(9618);
    outputs(2112) <= (layer2_outputs(8227)) or (layer2_outputs(533));
    outputs(2113) <= layer2_outputs(3915);
    outputs(2114) <= not(layer2_outputs(6515));
    outputs(2115) <= layer2_outputs(865);
    outputs(2116) <= (layer2_outputs(9952)) and not (layer2_outputs(301));
    outputs(2117) <= (layer2_outputs(2915)) xor (layer2_outputs(1863));
    outputs(2118) <= not((layer2_outputs(2880)) and (layer2_outputs(5253)));
    outputs(2119) <= layer2_outputs(6505);
    outputs(2120) <= not(layer2_outputs(2318));
    outputs(2121) <= not(layer2_outputs(4969));
    outputs(2122) <= layer2_outputs(3585);
    outputs(2123) <= not((layer2_outputs(4370)) and (layer2_outputs(6962)));
    outputs(2124) <= not(layer2_outputs(9633));
    outputs(2125) <= layer2_outputs(1714);
    outputs(2126) <= not(layer2_outputs(3146));
    outputs(2127) <= not(layer2_outputs(6353));
    outputs(2128) <= layer2_outputs(3272);
    outputs(2129) <= layer2_outputs(7585);
    outputs(2130) <= (layer2_outputs(1917)) or (layer2_outputs(9365));
    outputs(2131) <= (layer2_outputs(5635)) and not (layer2_outputs(9702));
    outputs(2132) <= (layer2_outputs(5013)) xor (layer2_outputs(6200));
    outputs(2133) <= not((layer2_outputs(2839)) xor (layer2_outputs(1107)));
    outputs(2134) <= (layer2_outputs(2913)) and not (layer2_outputs(1000));
    outputs(2135) <= not(layer2_outputs(290));
    outputs(2136) <= layer2_outputs(7596);
    outputs(2137) <= not((layer2_outputs(8768)) and (layer2_outputs(3041)));
    outputs(2138) <= layer2_outputs(6916);
    outputs(2139) <= (layer2_outputs(2871)) and (layer2_outputs(7469));
    outputs(2140) <= (layer2_outputs(231)) xor (layer2_outputs(9280));
    outputs(2141) <= layer2_outputs(3968);
    outputs(2142) <= not(layer2_outputs(1542));
    outputs(2143) <= not(layer2_outputs(9517));
    outputs(2144) <= layer2_outputs(3351);
    outputs(2145) <= not(layer2_outputs(7793));
    outputs(2146) <= not(layer2_outputs(726)) or (layer2_outputs(4564));
    outputs(2147) <= (layer2_outputs(3071)) xor (layer2_outputs(6320));
    outputs(2148) <= not((layer2_outputs(8577)) xor (layer2_outputs(2415)));
    outputs(2149) <= layer2_outputs(3840);
    outputs(2150) <= (layer2_outputs(8220)) or (layer2_outputs(6097));
    outputs(2151) <= not(layer2_outputs(923)) or (layer2_outputs(3438));
    outputs(2152) <= layer2_outputs(2632);
    outputs(2153) <= not(layer2_outputs(4346));
    outputs(2154) <= not(layer2_outputs(916));
    outputs(2155) <= not(layer2_outputs(3525));
    outputs(2156) <= not((layer2_outputs(6577)) xor (layer2_outputs(1737)));
    outputs(2157) <= (layer2_outputs(7986)) xor (layer2_outputs(1795));
    outputs(2158) <= not((layer2_outputs(3503)) xor (layer2_outputs(8569)));
    outputs(2159) <= layer2_outputs(8887);
    outputs(2160) <= (layer2_outputs(5074)) xor (layer2_outputs(4155));
    outputs(2161) <= (layer2_outputs(1914)) and (layer2_outputs(9398));
    outputs(2162) <= layer2_outputs(6669);
    outputs(2163) <= not(layer2_outputs(2881));
    outputs(2164) <= not(layer2_outputs(992)) or (layer2_outputs(7027));
    outputs(2165) <= not(layer2_outputs(7487));
    outputs(2166) <= layer2_outputs(2117);
    outputs(2167) <= (layer2_outputs(9968)) and not (layer2_outputs(2958));
    outputs(2168) <= not(layer2_outputs(6595));
    outputs(2169) <= not(layer2_outputs(2335));
    outputs(2170) <= layer2_outputs(8685);
    outputs(2171) <= not(layer2_outputs(8499));
    outputs(2172) <= not(layer2_outputs(7784));
    outputs(2173) <= (layer2_outputs(1109)) or (layer2_outputs(5013));
    outputs(2174) <= not(layer2_outputs(4425));
    outputs(2175) <= (layer2_outputs(10027)) and (layer2_outputs(5651));
    outputs(2176) <= layer2_outputs(4025);
    outputs(2177) <= not(layer2_outputs(660));
    outputs(2178) <= layer2_outputs(8516);
    outputs(2179) <= (layer2_outputs(2170)) xor (layer2_outputs(9229));
    outputs(2180) <= layer2_outputs(1889);
    outputs(2181) <= not(layer2_outputs(8706));
    outputs(2182) <= (layer2_outputs(2879)) or (layer2_outputs(3401));
    outputs(2183) <= not(layer2_outputs(6895));
    outputs(2184) <= layer2_outputs(4255);
    outputs(2185) <= not((layer2_outputs(5109)) and (layer2_outputs(9890)));
    outputs(2186) <= layer2_outputs(9467);
    outputs(2187) <= not(layer2_outputs(8689)) or (layer2_outputs(2304));
    outputs(2188) <= not(layer2_outputs(256));
    outputs(2189) <= not(layer2_outputs(7073));
    outputs(2190) <= layer2_outputs(8209);
    outputs(2191) <= not((layer2_outputs(2316)) xor (layer2_outputs(904)));
    outputs(2192) <= layer2_outputs(10196);
    outputs(2193) <= (layer2_outputs(10001)) xor (layer2_outputs(9869));
    outputs(2194) <= not(layer2_outputs(6278));
    outputs(2195) <= not((layer2_outputs(7715)) and (layer2_outputs(213)));
    outputs(2196) <= (layer2_outputs(10032)) and not (layer2_outputs(5907));
    outputs(2197) <= not(layer2_outputs(3347));
    outputs(2198) <= layer2_outputs(788);
    outputs(2199) <= not(layer2_outputs(4554));
    outputs(2200) <= not(layer2_outputs(1348)) or (layer2_outputs(3362));
    outputs(2201) <= (layer2_outputs(7848)) or (layer2_outputs(7217));
    outputs(2202) <= not(layer2_outputs(5737));
    outputs(2203) <= not(layer2_outputs(4743));
    outputs(2204) <= layer2_outputs(8524);
    outputs(2205) <= (layer2_outputs(3725)) or (layer2_outputs(10033));
    outputs(2206) <= (layer2_outputs(1870)) xor (layer2_outputs(9526));
    outputs(2207) <= layer2_outputs(6955);
    outputs(2208) <= not(layer2_outputs(19)) or (layer2_outputs(10074));
    outputs(2209) <= (layer2_outputs(3425)) xor (layer2_outputs(1373));
    outputs(2210) <= not((layer2_outputs(4287)) xor (layer2_outputs(8469)));
    outputs(2211) <= not(layer2_outputs(776)) or (layer2_outputs(5997));
    outputs(2212) <= not(layer2_outputs(1416)) or (layer2_outputs(7069));
    outputs(2213) <= layer2_outputs(10033);
    outputs(2214) <= (layer2_outputs(7014)) and not (layer2_outputs(291));
    outputs(2215) <= layer2_outputs(343);
    outputs(2216) <= layer2_outputs(3442);
    outputs(2217) <= (layer2_outputs(1754)) xor (layer2_outputs(2642));
    outputs(2218) <= layer2_outputs(3290);
    outputs(2219) <= layer2_outputs(7796);
    outputs(2220) <= (layer2_outputs(4605)) xor (layer2_outputs(8313));
    outputs(2221) <= layer2_outputs(3267);
    outputs(2222) <= not(layer2_outputs(8922));
    outputs(2223) <= (layer2_outputs(7614)) xor (layer2_outputs(9630));
    outputs(2224) <= (layer2_outputs(7963)) and not (layer2_outputs(7590));
    outputs(2225) <= (layer2_outputs(6869)) and (layer2_outputs(7882));
    outputs(2226) <= not((layer2_outputs(6708)) and (layer2_outputs(9757)));
    outputs(2227) <= not(layer2_outputs(5653)) or (layer2_outputs(1673));
    outputs(2228) <= not(layer2_outputs(9235));
    outputs(2229) <= layer2_outputs(5274);
    outputs(2230) <= layer2_outputs(5342);
    outputs(2231) <= not((layer2_outputs(6078)) xor (layer2_outputs(4005)));
    outputs(2232) <= layer2_outputs(9798);
    outputs(2233) <= (layer2_outputs(3804)) and (layer2_outputs(5224));
    outputs(2234) <= not(layer2_outputs(3256)) or (layer2_outputs(4998));
    outputs(2235) <= layer2_outputs(1236);
    outputs(2236) <= not(layer2_outputs(9060));
    outputs(2237) <= not(layer2_outputs(3984));
    outputs(2238) <= not((layer2_outputs(1941)) xor (layer2_outputs(3833)));
    outputs(2239) <= layer2_outputs(7121);
    outputs(2240) <= not(layer2_outputs(9464));
    outputs(2241) <= (layer2_outputs(7789)) xor (layer2_outputs(6427));
    outputs(2242) <= layer2_outputs(4062);
    outputs(2243) <= not(layer2_outputs(1975));
    outputs(2244) <= layer2_outputs(3986);
    outputs(2245) <= layer2_outputs(5536);
    outputs(2246) <= not((layer2_outputs(3031)) and (layer2_outputs(798)));
    outputs(2247) <= layer2_outputs(6745);
    outputs(2248) <= layer2_outputs(2586);
    outputs(2249) <= (layer2_outputs(1396)) and not (layer2_outputs(5120));
    outputs(2250) <= layer2_outputs(9272);
    outputs(2251) <= (layer2_outputs(3828)) and not (layer2_outputs(4746));
    outputs(2252) <= layer2_outputs(9140);
    outputs(2253) <= not((layer2_outputs(2277)) or (layer2_outputs(1396)));
    outputs(2254) <= not(layer2_outputs(4131));
    outputs(2255) <= not(layer2_outputs(5295));
    outputs(2256) <= (layer2_outputs(3978)) xor (layer2_outputs(1678));
    outputs(2257) <= not(layer2_outputs(8246));
    outputs(2258) <= layer2_outputs(9759);
    outputs(2259) <= not(layer2_outputs(3768));
    outputs(2260) <= (layer2_outputs(5888)) or (layer2_outputs(10153));
    outputs(2261) <= (layer2_outputs(6099)) xor (layer2_outputs(9640));
    outputs(2262) <= layer2_outputs(9777);
    outputs(2263) <= (layer2_outputs(1916)) or (layer2_outputs(6683));
    outputs(2264) <= not(layer2_outputs(4857));
    outputs(2265) <= not(layer2_outputs(552));
    outputs(2266) <= layer2_outputs(4732);
    outputs(2267) <= (layer2_outputs(5624)) or (layer2_outputs(4202));
    outputs(2268) <= (layer2_outputs(8189)) and not (layer2_outputs(3312));
    outputs(2269) <= not(layer2_outputs(9306));
    outputs(2270) <= layer2_outputs(7835);
    outputs(2271) <= not(layer2_outputs(9757)) or (layer2_outputs(2180));
    outputs(2272) <= not(layer2_outputs(9060));
    outputs(2273) <= layer2_outputs(10192);
    outputs(2274) <= not((layer2_outputs(3943)) and (layer2_outputs(3757)));
    outputs(2275) <= (layer2_outputs(7867)) and not (layer2_outputs(7942));
    outputs(2276) <= layer2_outputs(4299);
    outputs(2277) <= not(layer2_outputs(6026));
    outputs(2278) <= not((layer2_outputs(1558)) and (layer2_outputs(8886)));
    outputs(2279) <= not(layer2_outputs(1698));
    outputs(2280) <= not(layer2_outputs(9855));
    outputs(2281) <= not(layer2_outputs(4628));
    outputs(2282) <= not(layer2_outputs(4464)) or (layer2_outputs(2353));
    outputs(2283) <= (layer2_outputs(3731)) xor (layer2_outputs(749));
    outputs(2284) <= layer2_outputs(9883);
    outputs(2285) <= not(layer2_outputs(4109));
    outputs(2286) <= (layer2_outputs(281)) xor (layer2_outputs(10142));
    outputs(2287) <= layer2_outputs(1533);
    outputs(2288) <= not(layer2_outputs(7043));
    outputs(2289) <= not(layer2_outputs(7098));
    outputs(2290) <= layer2_outputs(9749);
    outputs(2291) <= layer2_outputs(932);
    outputs(2292) <= layer2_outputs(1581);
    outputs(2293) <= layer2_outputs(890);
    outputs(2294) <= not(layer2_outputs(6518)) or (layer2_outputs(4147));
    outputs(2295) <= layer2_outputs(2389);
    outputs(2296) <= not((layer2_outputs(4645)) or (layer2_outputs(4818)));
    outputs(2297) <= not((layer2_outputs(1241)) xor (layer2_outputs(8590)));
    outputs(2298) <= not((layer2_outputs(8419)) xor (layer2_outputs(6865)));
    outputs(2299) <= layer2_outputs(6839);
    outputs(2300) <= layer2_outputs(9087);
    outputs(2301) <= layer2_outputs(8807);
    outputs(2302) <= not((layer2_outputs(4174)) or (layer2_outputs(10190)));
    outputs(2303) <= (layer2_outputs(6633)) and (layer2_outputs(7064));
    outputs(2304) <= not((layer2_outputs(9416)) xor (layer2_outputs(6092)));
    outputs(2305) <= not(layer2_outputs(8307));
    outputs(2306) <= (layer2_outputs(9279)) xor (layer2_outputs(8386));
    outputs(2307) <= not(layer2_outputs(10219));
    outputs(2308) <= layer2_outputs(424);
    outputs(2309) <= layer2_outputs(5819);
    outputs(2310) <= (layer2_outputs(9912)) or (layer2_outputs(6910));
    outputs(2311) <= not((layer2_outputs(6488)) xor (layer2_outputs(382)));
    outputs(2312) <= layer2_outputs(3215);
    outputs(2313) <= layer2_outputs(2179);
    outputs(2314) <= (layer2_outputs(3687)) xor (layer2_outputs(7525));
    outputs(2315) <= layer2_outputs(9796);
    outputs(2316) <= layer2_outputs(1153);
    outputs(2317) <= layer2_outputs(5527);
    outputs(2318) <= (layer2_outputs(3741)) and not (layer2_outputs(7079));
    outputs(2319) <= (layer2_outputs(1543)) and (layer2_outputs(3571));
    outputs(2320) <= not(layer2_outputs(6984));
    outputs(2321) <= not(layer2_outputs(9075));
    outputs(2322) <= not((layer2_outputs(7905)) or (layer2_outputs(3375)));
    outputs(2323) <= not((layer2_outputs(7730)) or (layer2_outputs(8508)));
    outputs(2324) <= not(layer2_outputs(5994));
    outputs(2325) <= (layer2_outputs(3701)) xor (layer2_outputs(6240));
    outputs(2326) <= not(layer2_outputs(7201));
    outputs(2327) <= (layer2_outputs(3049)) xor (layer2_outputs(4682));
    outputs(2328) <= (layer2_outputs(725)) and (layer2_outputs(7750));
    outputs(2329) <= layer2_outputs(6433);
    outputs(2330) <= (layer2_outputs(8757)) and (layer2_outputs(1248));
    outputs(2331) <= (layer2_outputs(2874)) and (layer2_outputs(8197));
    outputs(2332) <= not(layer2_outputs(10194));
    outputs(2333) <= layer2_outputs(5186);
    outputs(2334) <= layer2_outputs(7585);
    outputs(2335) <= not(layer2_outputs(9659));
    outputs(2336) <= (layer2_outputs(10091)) xor (layer2_outputs(700));
    outputs(2337) <= (layer2_outputs(5643)) or (layer2_outputs(2252));
    outputs(2338) <= not(layer2_outputs(10133));
    outputs(2339) <= not((layer2_outputs(5511)) or (layer2_outputs(9205)));
    outputs(2340) <= layer2_outputs(7296);
    outputs(2341) <= not(layer2_outputs(3721));
    outputs(2342) <= (layer2_outputs(7341)) xor (layer2_outputs(1928));
    outputs(2343) <= not(layer2_outputs(9679));
    outputs(2344) <= not(layer2_outputs(7854)) or (layer2_outputs(4202));
    outputs(2345) <= layer2_outputs(8154);
    outputs(2346) <= layer2_outputs(8200);
    outputs(2347) <= not((layer2_outputs(5525)) xor (layer2_outputs(3131)));
    outputs(2348) <= layer2_outputs(79);
    outputs(2349) <= layer2_outputs(6448);
    outputs(2350) <= not(layer2_outputs(3213)) or (layer2_outputs(1955));
    outputs(2351) <= (layer2_outputs(3582)) and (layer2_outputs(8975));
    outputs(2352) <= not(layer2_outputs(6397));
    outputs(2353) <= not((layer2_outputs(2193)) or (layer2_outputs(2869)));
    outputs(2354) <= not((layer2_outputs(7009)) xor (layer2_outputs(8106)));
    outputs(2355) <= not(layer2_outputs(3563));
    outputs(2356) <= not(layer2_outputs(2334));
    outputs(2357) <= (layer2_outputs(4477)) xor (layer2_outputs(7621));
    outputs(2358) <= not((layer2_outputs(3906)) xor (layer2_outputs(6808)));
    outputs(2359) <= (layer2_outputs(2915)) and not (layer2_outputs(9762));
    outputs(2360) <= not(layer2_outputs(428));
    outputs(2361) <= not(layer2_outputs(6291));
    outputs(2362) <= layer2_outputs(6745);
    outputs(2363) <= layer2_outputs(1285);
    outputs(2364) <= (layer2_outputs(697)) and not (layer2_outputs(2384));
    outputs(2365) <= layer2_outputs(9516);
    outputs(2366) <= (layer2_outputs(3784)) and (layer2_outputs(586));
    outputs(2367) <= not(layer2_outputs(1157));
    outputs(2368) <= layer2_outputs(2709);
    outputs(2369) <= not(layer2_outputs(9053)) or (layer2_outputs(10107));
    outputs(2370) <= layer2_outputs(6920);
    outputs(2371) <= layer2_outputs(9525);
    outputs(2372) <= (layer2_outputs(796)) xor (layer2_outputs(2714));
    outputs(2373) <= layer2_outputs(2378);
    outputs(2374) <= not(layer2_outputs(7253));
    outputs(2375) <= not(layer2_outputs(572));
    outputs(2376) <= (layer2_outputs(4324)) or (layer2_outputs(7471));
    outputs(2377) <= layer2_outputs(5449);
    outputs(2378) <= (layer2_outputs(7858)) and (layer2_outputs(1183));
    outputs(2379) <= not(layer2_outputs(4594));
    outputs(2380) <= not(layer2_outputs(1160));
    outputs(2381) <= (layer2_outputs(2037)) xor (layer2_outputs(9651));
    outputs(2382) <= layer2_outputs(8348);
    outputs(2383) <= not(layer2_outputs(2490));
    outputs(2384) <= not((layer2_outputs(4894)) or (layer2_outputs(5514)));
    outputs(2385) <= layer2_outputs(3395);
    outputs(2386) <= (layer2_outputs(1696)) or (layer2_outputs(5398));
    outputs(2387) <= layer2_outputs(8645);
    outputs(2388) <= not(layer2_outputs(7397));
    outputs(2389) <= not(layer2_outputs(4033));
    outputs(2390) <= not(layer2_outputs(7534));
    outputs(2391) <= not((layer2_outputs(5169)) xor (layer2_outputs(1252)));
    outputs(2392) <= not(layer2_outputs(881)) or (layer2_outputs(5588));
    outputs(2393) <= (layer2_outputs(9842)) or (layer2_outputs(8853));
    outputs(2394) <= (layer2_outputs(9027)) and (layer2_outputs(2053));
    outputs(2395) <= not((layer2_outputs(6885)) xor (layer2_outputs(4900)));
    outputs(2396) <= not((layer2_outputs(2016)) xor (layer2_outputs(2865)));
    outputs(2397) <= not((layer2_outputs(1983)) or (layer2_outputs(7072)));
    outputs(2398) <= (layer2_outputs(8403)) xor (layer2_outputs(1731));
    outputs(2399) <= layer2_outputs(4485);
    outputs(2400) <= not(layer2_outputs(3572));
    outputs(2401) <= not(layer2_outputs(2730)) or (layer2_outputs(6489));
    outputs(2402) <= (layer2_outputs(2626)) and not (layer2_outputs(4472));
    outputs(2403) <= (layer2_outputs(4383)) xor (layer2_outputs(9007));
    outputs(2404) <= layer2_outputs(1488);
    outputs(2405) <= not((layer2_outputs(7812)) and (layer2_outputs(4710)));
    outputs(2406) <= not(layer2_outputs(319));
    outputs(2407) <= layer2_outputs(280);
    outputs(2408) <= (layer2_outputs(2536)) or (layer2_outputs(3544));
    outputs(2409) <= layer2_outputs(306);
    outputs(2410) <= not(layer2_outputs(4071)) or (layer2_outputs(1362));
    outputs(2411) <= (layer2_outputs(8104)) xor (layer2_outputs(7640));
    outputs(2412) <= layer2_outputs(3383);
    outputs(2413) <= not(layer2_outputs(10043));
    outputs(2414) <= (layer2_outputs(690)) and not (layer2_outputs(2243));
    outputs(2415) <= not(layer2_outputs(6392)) or (layer2_outputs(9244));
    outputs(2416) <= layer2_outputs(4130);
    outputs(2417) <= layer2_outputs(9131);
    outputs(2418) <= (layer2_outputs(5766)) and not (layer2_outputs(4520));
    outputs(2419) <= layer2_outputs(4558);
    outputs(2420) <= not(layer2_outputs(3643));
    outputs(2421) <= not(layer2_outputs(9740));
    outputs(2422) <= not(layer2_outputs(4916));
    outputs(2423) <= not((layer2_outputs(7236)) and (layer2_outputs(6932)));
    outputs(2424) <= not(layer2_outputs(6045));
    outputs(2425) <= not(layer2_outputs(3921));
    outputs(2426) <= not((layer2_outputs(9267)) or (layer2_outputs(1332)));
    outputs(2427) <= not(layer2_outputs(1347)) or (layer2_outputs(6830));
    outputs(2428) <= not(layer2_outputs(6715)) or (layer2_outputs(7599));
    outputs(2429) <= (layer2_outputs(5326)) or (layer2_outputs(2035));
    outputs(2430) <= layer2_outputs(935);
    outputs(2431) <= not(layer2_outputs(1399));
    outputs(2432) <= not(layer2_outputs(5814));
    outputs(2433) <= layer2_outputs(5354);
    outputs(2434) <= (layer2_outputs(5011)) and not (layer2_outputs(887));
    outputs(2435) <= not(layer2_outputs(7330));
    outputs(2436) <= not((layer2_outputs(7606)) xor (layer2_outputs(6142)));
    outputs(2437) <= layer2_outputs(7141);
    outputs(2438) <= not((layer2_outputs(3867)) xor (layer2_outputs(7108)));
    outputs(2439) <= layer2_outputs(7576);
    outputs(2440) <= not(layer2_outputs(1353)) or (layer2_outputs(3269));
    outputs(2441) <= not((layer2_outputs(9438)) xor (layer2_outputs(2867)));
    outputs(2442) <= not(layer2_outputs(866));
    outputs(2443) <= layer2_outputs(8378);
    outputs(2444) <= not(layer2_outputs(278));
    outputs(2445) <= layer2_outputs(4221);
    outputs(2446) <= not((layer2_outputs(3237)) xor (layer2_outputs(734)));
    outputs(2447) <= not(layer2_outputs(1613));
    outputs(2448) <= not(layer2_outputs(2497));
    outputs(2449) <= (layer2_outputs(5244)) xor (layer2_outputs(6924));
    outputs(2450) <= not(layer2_outputs(4550));
    outputs(2451) <= not(layer2_outputs(7365));
    outputs(2452) <= not(layer2_outputs(216)) or (layer2_outputs(2584));
    outputs(2453) <= not((layer2_outputs(9440)) xor (layer2_outputs(5883)));
    outputs(2454) <= not(layer2_outputs(1124));
    outputs(2455) <= (layer2_outputs(2094)) xor (layer2_outputs(10040));
    outputs(2456) <= not(layer2_outputs(8957)) or (layer2_outputs(6611));
    outputs(2457) <= not(layer2_outputs(3113)) or (layer2_outputs(8033));
    outputs(2458) <= layer2_outputs(1583);
    outputs(2459) <= (layer2_outputs(6058)) xor (layer2_outputs(3405));
    outputs(2460) <= not(layer2_outputs(8185));
    outputs(2461) <= not(layer2_outputs(3042));
    outputs(2462) <= (layer2_outputs(8208)) or (layer2_outputs(7822));
    outputs(2463) <= layer2_outputs(5418);
    outputs(2464) <= not((layer2_outputs(9542)) or (layer2_outputs(6099)));
    outputs(2465) <= not(layer2_outputs(8545));
    outputs(2466) <= layer2_outputs(4235);
    outputs(2467) <= layer2_outputs(4427);
    outputs(2468) <= not(layer2_outputs(204));
    outputs(2469) <= not(layer2_outputs(9710));
    outputs(2470) <= (layer2_outputs(4120)) and not (layer2_outputs(1895));
    outputs(2471) <= not((layer2_outputs(6782)) and (layer2_outputs(9795)));
    outputs(2472) <= layer2_outputs(2676);
    outputs(2473) <= not(layer2_outputs(4055)) or (layer2_outputs(311));
    outputs(2474) <= not(layer2_outputs(2652));
    outputs(2475) <= not((layer2_outputs(1796)) and (layer2_outputs(3875)));
    outputs(2476) <= not((layer2_outputs(1197)) xor (layer2_outputs(2171)));
    outputs(2477) <= (layer2_outputs(9171)) xor (layer2_outputs(3552));
    outputs(2478) <= not((layer2_outputs(9566)) xor (layer2_outputs(2622)));
    outputs(2479) <= layer2_outputs(703);
    outputs(2480) <= layer2_outputs(9005);
    outputs(2481) <= layer2_outputs(5390);
    outputs(2482) <= layer2_outputs(6046);
    outputs(2483) <= not(layer2_outputs(6723)) or (layer2_outputs(5618));
    outputs(2484) <= not((layer2_outputs(8317)) xor (layer2_outputs(1929)));
    outputs(2485) <= not(layer2_outputs(2065));
    outputs(2486) <= layer2_outputs(431);
    outputs(2487) <= (layer2_outputs(6645)) xor (layer2_outputs(7262));
    outputs(2488) <= not(layer2_outputs(2250));
    outputs(2489) <= layer2_outputs(2571);
    outputs(2490) <= layer2_outputs(8623);
    outputs(2491) <= not(layer2_outputs(1124));
    outputs(2492) <= layer2_outputs(4208);
    outputs(2493) <= layer2_outputs(2638);
    outputs(2494) <= not(layer2_outputs(3143));
    outputs(2495) <= (layer2_outputs(2274)) and (layer2_outputs(1359));
    outputs(2496) <= not(layer2_outputs(1608));
    outputs(2497) <= not(layer2_outputs(1622));
    outputs(2498) <= layer2_outputs(6572);
    outputs(2499) <= layer2_outputs(996);
    outputs(2500) <= layer2_outputs(3691);
    outputs(2501) <= not(layer2_outputs(364));
    outputs(2502) <= (layer2_outputs(10068)) xor (layer2_outputs(987));
    outputs(2503) <= not(layer2_outputs(5587));
    outputs(2504) <= layer2_outputs(9806);
    outputs(2505) <= not(layer2_outputs(9578));
    outputs(2506) <= not(layer2_outputs(2559));
    outputs(2507) <= layer2_outputs(8043);
    outputs(2508) <= not(layer2_outputs(7144));
    outputs(2509) <= (layer2_outputs(9305)) or (layer2_outputs(7492));
    outputs(2510) <= layer2_outputs(1049);
    outputs(2511) <= layer2_outputs(6083);
    outputs(2512) <= not((layer2_outputs(9352)) xor (layer2_outputs(5243)));
    outputs(2513) <= (layer2_outputs(9981)) or (layer2_outputs(2026));
    outputs(2514) <= layer2_outputs(3777);
    outputs(2515) <= not(layer2_outputs(6091));
    outputs(2516) <= (layer2_outputs(1744)) xor (layer2_outputs(6912));
    outputs(2517) <= not(layer2_outputs(6339));
    outputs(2518) <= layer2_outputs(2376);
    outputs(2519) <= not(layer2_outputs(8055));
    outputs(2520) <= (layer2_outputs(29)) xor (layer2_outputs(8738));
    outputs(2521) <= layer2_outputs(2097);
    outputs(2522) <= not((layer2_outputs(1424)) or (layer2_outputs(8291)));
    outputs(2523) <= layer2_outputs(484);
    outputs(2524) <= not(layer2_outputs(9354)) or (layer2_outputs(9751));
    outputs(2525) <= layer2_outputs(802);
    outputs(2526) <= layer2_outputs(1383);
    outputs(2527) <= not((layer2_outputs(3966)) and (layer2_outputs(1477)));
    outputs(2528) <= not(layer2_outputs(1768));
    outputs(2529) <= (layer2_outputs(419)) and not (layer2_outputs(2321));
    outputs(2530) <= layer2_outputs(9706);
    outputs(2531) <= (layer2_outputs(9609)) xor (layer2_outputs(1048));
    outputs(2532) <= (layer2_outputs(6288)) and (layer2_outputs(8576));
    outputs(2533) <= not(layer2_outputs(551));
    outputs(2534) <= layer2_outputs(78);
    outputs(2535) <= not(layer2_outputs(1060));
    outputs(2536) <= (layer2_outputs(4104)) and not (layer2_outputs(6159));
    outputs(2537) <= (layer2_outputs(870)) xor (layer2_outputs(8953));
    outputs(2538) <= layer2_outputs(2133);
    outputs(2539) <= (layer2_outputs(37)) xor (layer2_outputs(8311));
    outputs(2540) <= not(layer2_outputs(4304)) or (layer2_outputs(1024));
    outputs(2541) <= (layer2_outputs(9766)) and not (layer2_outputs(9158));
    outputs(2542) <= not(layer2_outputs(2084));
    outputs(2543) <= layer2_outputs(3849);
    outputs(2544) <= not(layer2_outputs(6546));
    outputs(2545) <= not(layer2_outputs(4007));
    outputs(2546) <= not(layer2_outputs(9170));
    outputs(2547) <= not(layer2_outputs(9003));
    outputs(2548) <= (layer2_outputs(6926)) or (layer2_outputs(3184));
    outputs(2549) <= not(layer2_outputs(6407));
    outputs(2550) <= layer2_outputs(4578);
    outputs(2551) <= not(layer2_outputs(2653));
    outputs(2552) <= (layer2_outputs(4882)) and not (layer2_outputs(1937));
    outputs(2553) <= not(layer2_outputs(6026));
    outputs(2554) <= not((layer2_outputs(9578)) or (layer2_outputs(10085)));
    outputs(2555) <= not(layer2_outputs(2410));
    outputs(2556) <= not((layer2_outputs(7875)) and (layer2_outputs(2282)));
    outputs(2557) <= (layer2_outputs(627)) or (layer2_outputs(2493));
    outputs(2558) <= layer2_outputs(4591);
    outputs(2559) <= layer2_outputs(8416);
    outputs(2560) <= not(layer2_outputs(6617)) or (layer2_outputs(3184));
    outputs(2561) <= not(layer2_outputs(6804));
    outputs(2562) <= (layer2_outputs(2928)) xor (layer2_outputs(6249));
    outputs(2563) <= (layer2_outputs(7316)) xor (layer2_outputs(2663));
    outputs(2564) <= (layer2_outputs(373)) and not (layer2_outputs(847));
    outputs(2565) <= layer2_outputs(933);
    outputs(2566) <= not(layer2_outputs(4819));
    outputs(2567) <= not((layer2_outputs(8913)) and (layer2_outputs(8014)));
    outputs(2568) <= (layer2_outputs(4373)) xor (layer2_outputs(8727));
    outputs(2569) <= not((layer2_outputs(4783)) xor (layer2_outputs(19)));
    outputs(2570) <= not(layer2_outputs(7450));
    outputs(2571) <= layer2_outputs(4127);
    outputs(2572) <= layer2_outputs(8690);
    outputs(2573) <= not(layer2_outputs(1964));
    outputs(2574) <= layer2_outputs(3638);
    outputs(2575) <= not((layer2_outputs(7241)) xor (layer2_outputs(4034)));
    outputs(2576) <= layer2_outputs(3450);
    outputs(2577) <= not((layer2_outputs(6674)) or (layer2_outputs(8752)));
    outputs(2578) <= not(layer2_outputs(1384));
    outputs(2579) <= not((layer2_outputs(7739)) and (layer2_outputs(2045)));
    outputs(2580) <= not((layer2_outputs(5589)) xor (layer2_outputs(9720)));
    outputs(2581) <= not(layer2_outputs(8507));
    outputs(2582) <= layer2_outputs(7952);
    outputs(2583) <= not(layer2_outputs(7438));
    outputs(2584) <= not(layer2_outputs(9964));
    outputs(2585) <= layer2_outputs(5580);
    outputs(2586) <= layer2_outputs(8101);
    outputs(2587) <= not(layer2_outputs(8572));
    outputs(2588) <= not(layer2_outputs(9190));
    outputs(2589) <= layer2_outputs(8867);
    outputs(2590) <= (layer2_outputs(9945)) xor (layer2_outputs(1759));
    outputs(2591) <= not(layer2_outputs(316));
    outputs(2592) <= not(layer2_outputs(3103));
    outputs(2593) <= not((layer2_outputs(5191)) xor (layer2_outputs(4825)));
    outputs(2594) <= not(layer2_outputs(470));
    outputs(2595) <= not(layer2_outputs(9298));
    outputs(2596) <= not((layer2_outputs(4083)) xor (layer2_outputs(2710)));
    outputs(2597) <= not(layer2_outputs(4822)) or (layer2_outputs(10000));
    outputs(2598) <= (layer2_outputs(1397)) and (layer2_outputs(1511));
    outputs(2599) <= not(layer2_outputs(5871));
    outputs(2600) <= not(layer2_outputs(7387)) or (layer2_outputs(3971));
    outputs(2601) <= layer2_outputs(7468);
    outputs(2602) <= layer2_outputs(5757);
    outputs(2603) <= not(layer2_outputs(516));
    outputs(2604) <= not(layer2_outputs(9917));
    outputs(2605) <= not(layer2_outputs(4343));
    outputs(2606) <= not((layer2_outputs(215)) xor (layer2_outputs(6602)));
    outputs(2607) <= layer2_outputs(5921);
    outputs(2608) <= not(layer2_outputs(5693)) or (layer2_outputs(6655));
    outputs(2609) <= (layer2_outputs(4123)) and not (layer2_outputs(5886));
    outputs(2610) <= (layer2_outputs(5285)) and not (layer2_outputs(3729));
    outputs(2611) <= not(layer2_outputs(3945));
    outputs(2612) <= layer2_outputs(8249);
    outputs(2613) <= (layer2_outputs(3234)) or (layer2_outputs(1208));
    outputs(2614) <= layer2_outputs(10088);
    outputs(2615) <= not(layer2_outputs(7413));
    outputs(2616) <= not(layer2_outputs(8994));
    outputs(2617) <= not(layer2_outputs(901));
    outputs(2618) <= (layer2_outputs(5932)) or (layer2_outputs(6189));
    outputs(2619) <= (layer2_outputs(9313)) and not (layer2_outputs(383));
    outputs(2620) <= not(layer2_outputs(9044)) or (layer2_outputs(1741));
    outputs(2621) <= not(layer2_outputs(4556)) or (layer2_outputs(4154));
    outputs(2622) <= not(layer2_outputs(6210));
    outputs(2623) <= not(layer2_outputs(7345));
    outputs(2624) <= not(layer2_outputs(6835));
    outputs(2625) <= not((layer2_outputs(10160)) xor (layer2_outputs(6778)));
    outputs(2626) <= not((layer2_outputs(7887)) and (layer2_outputs(6583)));
    outputs(2627) <= layer2_outputs(8149);
    outputs(2628) <= not(layer2_outputs(7302));
    outputs(2629) <= layer2_outputs(1049);
    outputs(2630) <= layer2_outputs(3457);
    outputs(2631) <= not(layer2_outputs(8298)) or (layer2_outputs(8787));
    outputs(2632) <= not(layer2_outputs(5365));
    outputs(2633) <= (layer2_outputs(3869)) xor (layer2_outputs(2011));
    outputs(2634) <= layer2_outputs(5728);
    outputs(2635) <= not(layer2_outputs(3662));
    outputs(2636) <= not((layer2_outputs(10106)) xor (layer2_outputs(1538)));
    outputs(2637) <= not((layer2_outputs(73)) and (layer2_outputs(135)));
    outputs(2638) <= layer2_outputs(9736);
    outputs(2639) <= not((layer2_outputs(1999)) xor (layer2_outputs(450)));
    outputs(2640) <= layer2_outputs(3791);
    outputs(2641) <= (layer2_outputs(4502)) xor (layer2_outputs(5647));
    outputs(2642) <= layer2_outputs(3797);
    outputs(2643) <= not(layer2_outputs(6690));
    outputs(2644) <= layer2_outputs(3580);
    outputs(2645) <= layer2_outputs(511);
    outputs(2646) <= layer2_outputs(9087);
    outputs(2647) <= not((layer2_outputs(3348)) xor (layer2_outputs(6763)));
    outputs(2648) <= not((layer2_outputs(10148)) xor (layer2_outputs(5494)));
    outputs(2649) <= layer2_outputs(1027);
    outputs(2650) <= not(layer2_outputs(4377));
    outputs(2651) <= not(layer2_outputs(1510));
    outputs(2652) <= not(layer2_outputs(4)) or (layer2_outputs(7310));
    outputs(2653) <= not(layer2_outputs(9182));
    outputs(2654) <= layer2_outputs(6181);
    outputs(2655) <= not(layer2_outputs(6272));
    outputs(2656) <= not(layer2_outputs(6283));
    outputs(2657) <= (layer2_outputs(6335)) and not (layer2_outputs(10172));
    outputs(2658) <= not(layer2_outputs(1080)) or (layer2_outputs(5681));
    outputs(2659) <= not((layer2_outputs(905)) xor (layer2_outputs(2048)));
    outputs(2660) <= layer2_outputs(3626);
    outputs(2661) <= not(layer2_outputs(1833));
    outputs(2662) <= layer2_outputs(6748);
    outputs(2663) <= not((layer2_outputs(432)) xor (layer2_outputs(9900)));
    outputs(2664) <= (layer2_outputs(6797)) and (layer2_outputs(367));
    outputs(2665) <= not(layer2_outputs(9404));
    outputs(2666) <= layer2_outputs(4162);
    outputs(2667) <= layer2_outputs(8339);
    outputs(2668) <= layer2_outputs(3794);
    outputs(2669) <= (layer2_outputs(2983)) and not (layer2_outputs(5736));
    outputs(2670) <= not(layer2_outputs(1229));
    outputs(2671) <= layer2_outputs(1350);
    outputs(2672) <= layer2_outputs(8843);
    outputs(2673) <= (layer2_outputs(4300)) xor (layer2_outputs(349));
    outputs(2674) <= layer2_outputs(9189);
    outputs(2675) <= layer2_outputs(8267);
    outputs(2676) <= not((layer2_outputs(2975)) xor (layer2_outputs(150)));
    outputs(2677) <= not(layer2_outputs(634));
    outputs(2678) <= layer2_outputs(2603);
    outputs(2679) <= (layer2_outputs(8902)) and not (layer2_outputs(4179));
    outputs(2680) <= (layer2_outputs(9178)) or (layer2_outputs(4271));
    outputs(2681) <= not(layer2_outputs(8919)) or (layer2_outputs(1299));
    outputs(2682) <= not((layer2_outputs(247)) xor (layer2_outputs(1936)));
    outputs(2683) <= (layer2_outputs(1600)) xor (layer2_outputs(7918));
    outputs(2684) <= layer2_outputs(5199);
    outputs(2685) <= layer2_outputs(6799);
    outputs(2686) <= layer2_outputs(8378);
    outputs(2687) <= (layer2_outputs(9073)) and not (layer2_outputs(7264));
    outputs(2688) <= (layer2_outputs(6142)) xor (layer2_outputs(1802));
    outputs(2689) <= (layer2_outputs(6952)) and not (layer2_outputs(6811));
    outputs(2690) <= not((layer2_outputs(5236)) xor (layer2_outputs(4843)));
    outputs(2691) <= not((layer2_outputs(1998)) xor (layer2_outputs(5629)));
    outputs(2692) <= not(layer2_outputs(1856)) or (layer2_outputs(147));
    outputs(2693) <= not(layer2_outputs(9012));
    outputs(2694) <= (layer2_outputs(5779)) and (layer2_outputs(7496));
    outputs(2695) <= layer2_outputs(420);
    outputs(2696) <= (layer2_outputs(6845)) and not (layer2_outputs(2433));
    outputs(2697) <= (layer2_outputs(10184)) and not (layer2_outputs(9810));
    outputs(2698) <= not(layer2_outputs(682));
    outputs(2699) <= not(layer2_outputs(7265));
    outputs(2700) <= not(layer2_outputs(9255));
    outputs(2701) <= layer2_outputs(303);
    outputs(2702) <= (layer2_outputs(5519)) and (layer2_outputs(3715));
    outputs(2703) <= layer2_outputs(5688);
    outputs(2704) <= not(layer2_outputs(6834));
    outputs(2705) <= layer2_outputs(6838);
    outputs(2706) <= not((layer2_outputs(8680)) xor (layer2_outputs(9992)));
    outputs(2707) <= not(layer2_outputs(6665));
    outputs(2708) <= not((layer2_outputs(1918)) xor (layer2_outputs(7303)));
    outputs(2709) <= (layer2_outputs(7691)) xor (layer2_outputs(1620));
    outputs(2710) <= not(layer2_outputs(2708)) or (layer2_outputs(8544));
    outputs(2711) <= not(layer2_outputs(9327));
    outputs(2712) <= not((layer2_outputs(6101)) and (layer2_outputs(3663)));
    outputs(2713) <= not((layer2_outputs(5158)) xor (layer2_outputs(6109)));
    outputs(2714) <= layer2_outputs(2409);
    outputs(2715) <= layer2_outputs(10083);
    outputs(2716) <= (layer2_outputs(714)) and not (layer2_outputs(9718));
    outputs(2717) <= '1';
    outputs(2718) <= (layer2_outputs(6987)) xor (layer2_outputs(8420));
    outputs(2719) <= not((layer2_outputs(9441)) xor (layer2_outputs(4078)));
    outputs(2720) <= layer2_outputs(6234);
    outputs(2721) <= not(layer2_outputs(3936)) or (layer2_outputs(10075));
    outputs(2722) <= layer2_outputs(9294);
    outputs(2723) <= layer2_outputs(6404);
    outputs(2724) <= (layer2_outputs(785)) or (layer2_outputs(8376));
    outputs(2725) <= layer2_outputs(5132);
    outputs(2726) <= layer2_outputs(1198);
    outputs(2727) <= not((layer2_outputs(9860)) or (layer2_outputs(8470)));
    outputs(2728) <= layer2_outputs(7852);
    outputs(2729) <= layer2_outputs(3445);
    outputs(2730) <= not(layer2_outputs(7327));
    outputs(2731) <= not(layer2_outputs(5487)) or (layer2_outputs(4084));
    outputs(2732) <= not(layer2_outputs(2964));
    outputs(2733) <= not(layer2_outputs(8764));
    outputs(2734) <= (layer2_outputs(2008)) xor (layer2_outputs(8415));
    outputs(2735) <= not((layer2_outputs(5984)) or (layer2_outputs(914)));
    outputs(2736) <= layer2_outputs(8753);
    outputs(2737) <= (layer2_outputs(902)) xor (layer2_outputs(8772));
    outputs(2738) <= layer2_outputs(184);
    outputs(2739) <= not(layer2_outputs(3672));
    outputs(2740) <= not((layer2_outputs(5577)) xor (layer2_outputs(1462)));
    outputs(2741) <= not((layer2_outputs(5000)) xor (layer2_outputs(8418)));
    outputs(2742) <= not(layer2_outputs(2424));
    outputs(2743) <= not(layer2_outputs(1229));
    outputs(2744) <= not(layer2_outputs(9291));
    outputs(2745) <= not(layer2_outputs(2112));
    outputs(2746) <= (layer2_outputs(9960)) xor (layer2_outputs(4811));
    outputs(2747) <= layer2_outputs(9098);
    outputs(2748) <= not((layer2_outputs(10143)) xor (layer2_outputs(2561)));
    outputs(2749) <= layer2_outputs(3380);
    outputs(2750) <= not(layer2_outputs(1607)) or (layer2_outputs(4877));
    outputs(2751) <= not(layer2_outputs(7178));
    outputs(2752) <= not(layer2_outputs(6030));
    outputs(2753) <= not(layer2_outputs(7444));
    outputs(2754) <= (layer2_outputs(1365)) xor (layer2_outputs(3164));
    outputs(2755) <= layer2_outputs(5850);
    outputs(2756) <= not((layer2_outputs(9788)) or (layer2_outputs(3618)));
    outputs(2757) <= layer2_outputs(5407);
    outputs(2758) <= (layer2_outputs(2123)) and (layer2_outputs(8286));
    outputs(2759) <= layer2_outputs(2666);
    outputs(2760) <= not(layer2_outputs(7707));
    outputs(2761) <= layer2_outputs(2404);
    outputs(2762) <= not(layer2_outputs(9125)) or (layer2_outputs(9240));
    outputs(2763) <= (layer2_outputs(1699)) or (layer2_outputs(8088));
    outputs(2764) <= layer2_outputs(2521);
    outputs(2765) <= layer2_outputs(137);
    outputs(2766) <= layer2_outputs(8702);
    outputs(2767) <= layer2_outputs(6188);
    outputs(2768) <= not(layer2_outputs(5509));
    outputs(2769) <= layer2_outputs(2977);
    outputs(2770) <= layer2_outputs(9513);
    outputs(2771) <= (layer2_outputs(4589)) or (layer2_outputs(6222));
    outputs(2772) <= not(layer2_outputs(219));
    outputs(2773) <= not(layer2_outputs(4990));
    outputs(2774) <= layer2_outputs(2153);
    outputs(2775) <= (layer2_outputs(4888)) xor (layer2_outputs(6054));
    outputs(2776) <= layer2_outputs(4030);
    outputs(2777) <= not(layer2_outputs(8147));
    outputs(2778) <= not((layer2_outputs(496)) xor (layer2_outputs(2640)));
    outputs(2779) <= not(layer2_outputs(7334));
    outputs(2780) <= not(layer2_outputs(8035));
    outputs(2781) <= layer2_outputs(5976);
    outputs(2782) <= layer2_outputs(8878);
    outputs(2783) <= (layer2_outputs(8654)) and not (layer2_outputs(9619));
    outputs(2784) <= (layer2_outputs(10156)) or (layer2_outputs(3744));
    outputs(2785) <= layer2_outputs(8180);
    outputs(2786) <= not((layer2_outputs(2083)) or (layer2_outputs(8139)));
    outputs(2787) <= layer2_outputs(2545);
    outputs(2788) <= layer2_outputs(722);
    outputs(2789) <= not((layer2_outputs(1326)) xor (layer2_outputs(7919)));
    outputs(2790) <= not(layer2_outputs(2890));
    outputs(2791) <= layer2_outputs(2527);
    outputs(2792) <= not(layer2_outputs(651));
    outputs(2793) <= (layer2_outputs(1609)) xor (layer2_outputs(2109));
    outputs(2794) <= not(layer2_outputs(7397));
    outputs(2795) <= (layer2_outputs(3393)) and not (layer2_outputs(6062));
    outputs(2796) <= not(layer2_outputs(2459));
    outputs(2797) <= not((layer2_outputs(2866)) xor (layer2_outputs(10163)));
    outputs(2798) <= not(layer2_outputs(7618));
    outputs(2799) <= not(layer2_outputs(7439));
    outputs(2800) <= layer2_outputs(5521);
    outputs(2801) <= layer2_outputs(5255);
    outputs(2802) <= not(layer2_outputs(9799));
    outputs(2803) <= not(layer2_outputs(9739)) or (layer2_outputs(7176));
    outputs(2804) <= not((layer2_outputs(3015)) and (layer2_outputs(5717)));
    outputs(2805) <= not(layer2_outputs(10219));
    outputs(2806) <= not(layer2_outputs(3559)) or (layer2_outputs(2784));
    outputs(2807) <= layer2_outputs(309);
    outputs(2808) <= (layer2_outputs(1805)) and not (layer2_outputs(1015));
    outputs(2809) <= layer2_outputs(4226);
    outputs(2810) <= (layer2_outputs(6621)) or (layer2_outputs(1339));
    outputs(2811) <= layer2_outputs(8881);
    outputs(2812) <= not(layer2_outputs(5295));
    outputs(2813) <= not(layer2_outputs(1436));
    outputs(2814) <= not((layer2_outputs(6017)) xor (layer2_outputs(2850)));
    outputs(2815) <= layer2_outputs(6911);
    outputs(2816) <= layer2_outputs(9500);
    outputs(2817) <= (layer2_outputs(815)) xor (layer2_outputs(2098));
    outputs(2818) <= layer2_outputs(234);
    outputs(2819) <= layer2_outputs(6710);
    outputs(2820) <= (layer2_outputs(1735)) and (layer2_outputs(6946));
    outputs(2821) <= (layer2_outputs(2803)) and not (layer2_outputs(10189));
    outputs(2822) <= not(layer2_outputs(1817));
    outputs(2823) <= not(layer2_outputs(425));
    outputs(2824) <= not(layer2_outputs(3333));
    outputs(2825) <= not(layer2_outputs(9498));
    outputs(2826) <= not(layer2_outputs(1168));
    outputs(2827) <= (layer2_outputs(5005)) and not (layer2_outputs(3762));
    outputs(2828) <= not(layer2_outputs(692));
    outputs(2829) <= not(layer2_outputs(5576));
    outputs(2830) <= (layer2_outputs(3596)) or (layer2_outputs(8229));
    outputs(2831) <= not((layer2_outputs(7445)) xor (layer2_outputs(6354)));
    outputs(2832) <= layer2_outputs(1114);
    outputs(2833) <= (layer2_outputs(1032)) xor (layer2_outputs(1074));
    outputs(2834) <= not(layer2_outputs(8360));
    outputs(2835) <= not(layer2_outputs(1596)) or (layer2_outputs(528));
    outputs(2836) <= not(layer2_outputs(3444)) or (layer2_outputs(8571));
    outputs(2837) <= (layer2_outputs(9446)) xor (layer2_outputs(763));
    outputs(2838) <= not((layer2_outputs(10177)) xor (layer2_outputs(5444)));
    outputs(2839) <= layer2_outputs(8625);
    outputs(2840) <= layer2_outputs(151);
    outputs(2841) <= layer2_outputs(10169);
    outputs(2842) <= not((layer2_outputs(2906)) or (layer2_outputs(3497)));
    outputs(2843) <= layer2_outputs(1791);
    outputs(2844) <= not(layer2_outputs(2096));
    outputs(2845) <= not(layer2_outputs(122)) or (layer2_outputs(601));
    outputs(2846) <= not(layer2_outputs(4091));
    outputs(2847) <= layer2_outputs(890);
    outputs(2848) <= not((layer2_outputs(7893)) or (layer2_outputs(6242)));
    outputs(2849) <= layer2_outputs(1106);
    outputs(2850) <= not(layer2_outputs(794));
    outputs(2851) <= not(layer2_outputs(1896));
    outputs(2852) <= (layer2_outputs(6965)) and not (layer2_outputs(3757));
    outputs(2853) <= not(layer2_outputs(6201));
    outputs(2854) <= (layer2_outputs(7442)) xor (layer2_outputs(2416));
    outputs(2855) <= not((layer2_outputs(3963)) and (layer2_outputs(783)));
    outputs(2856) <= (layer2_outputs(8423)) and not (layer2_outputs(4327));
    outputs(2857) <= not(layer2_outputs(4832));
    outputs(2858) <= not(layer2_outputs(5730));
    outputs(2859) <= layer2_outputs(6308);
    outputs(2860) <= layer2_outputs(5445);
    outputs(2861) <= layer2_outputs(1183);
    outputs(2862) <= not(layer2_outputs(6549));
    outputs(2863) <= not(layer2_outputs(4270)) or (layer2_outputs(215));
    outputs(2864) <= layer2_outputs(6466);
    outputs(2865) <= layer2_outputs(7202);
    outputs(2866) <= not(layer2_outputs(2806)) or (layer2_outputs(7111));
    outputs(2867) <= not(layer2_outputs(5570));
    outputs(2868) <= layer2_outputs(10197);
    outputs(2869) <= not((layer2_outputs(5392)) xor (layer2_outputs(9870)));
    outputs(2870) <= (layer2_outputs(7866)) xor (layer2_outputs(647));
    outputs(2871) <= layer2_outputs(4622);
    outputs(2872) <= layer2_outputs(9593);
    outputs(2873) <= not((layer2_outputs(7385)) xor (layer2_outputs(8863)));
    outputs(2874) <= not((layer2_outputs(9580)) and (layer2_outputs(3719)));
    outputs(2875) <= (layer2_outputs(9136)) xor (layer2_outputs(2007));
    outputs(2876) <= (layer2_outputs(8211)) and not (layer2_outputs(3194));
    outputs(2877) <= not(layer2_outputs(348));
    outputs(2878) <= not((layer2_outputs(8943)) and (layer2_outputs(7995)));
    outputs(2879) <= not(layer2_outputs(1232));
    outputs(2880) <= layer2_outputs(258);
    outputs(2881) <= (layer2_outputs(7391)) xor (layer2_outputs(9020));
    outputs(2882) <= (layer2_outputs(7018)) and not (layer2_outputs(6087));
    outputs(2883) <= (layer2_outputs(3053)) xor (layer2_outputs(3404));
    outputs(2884) <= not((layer2_outputs(4640)) or (layer2_outputs(2616)));
    outputs(2885) <= not(layer2_outputs(1550));
    outputs(2886) <= not(layer2_outputs(4976));
    outputs(2887) <= not((layer2_outputs(1066)) xor (layer2_outputs(4426)));
    outputs(2888) <= layer2_outputs(8397);
    outputs(2889) <= not(layer2_outputs(422));
    outputs(2890) <= not(layer2_outputs(5737));
    outputs(2891) <= (layer2_outputs(6928)) or (layer2_outputs(1708));
    outputs(2892) <= (layer2_outputs(7409)) xor (layer2_outputs(4076));
    outputs(2893) <= (layer2_outputs(6937)) xor (layer2_outputs(9010));
    outputs(2894) <= layer2_outputs(4761);
    outputs(2895) <= (layer2_outputs(4230)) and not (layer2_outputs(2406));
    outputs(2896) <= (layer2_outputs(1295)) or (layer2_outputs(8153));
    outputs(2897) <= layer2_outputs(4000);
    outputs(2898) <= (layer2_outputs(2859)) and (layer2_outputs(3878));
    outputs(2899) <= layer2_outputs(9187);
    outputs(2900) <= layer2_outputs(6473);
    outputs(2901) <= not((layer2_outputs(9857)) xor (layer2_outputs(8999)));
    outputs(2902) <= (layer2_outputs(4111)) and (layer2_outputs(4974));
    outputs(2903) <= layer2_outputs(1592);
    outputs(2904) <= (layer2_outputs(3885)) xor (layer2_outputs(9518));
    outputs(2905) <= not(layer2_outputs(5113));
    outputs(2906) <= (layer2_outputs(6949)) or (layer2_outputs(6398));
    outputs(2907) <= (layer2_outputs(5332)) or (layer2_outputs(5479));
    outputs(2908) <= not(layer2_outputs(4587));
    outputs(2909) <= not(layer2_outputs(3931));
    outputs(2910) <= not(layer2_outputs(2290));
    outputs(2911) <= not(layer2_outputs(8330));
    outputs(2912) <= layer2_outputs(8175);
    outputs(2913) <= layer2_outputs(7939);
    outputs(2914) <= (layer2_outputs(7325)) xor (layer2_outputs(9219));
    outputs(2915) <= layer2_outputs(5313);
    outputs(2916) <= not(layer2_outputs(8167));
    outputs(2917) <= layer2_outputs(10167);
    outputs(2918) <= layer2_outputs(5789);
    outputs(2919) <= not(layer2_outputs(5423));
    outputs(2920) <= not(layer2_outputs(1953));
    outputs(2921) <= not(layer2_outputs(4641));
    outputs(2922) <= (layer2_outputs(7985)) and (layer2_outputs(6647));
    outputs(2923) <= not((layer2_outputs(5930)) xor (layer2_outputs(8018)));
    outputs(2924) <= not(layer2_outputs(7612));
    outputs(2925) <= not(layer2_outputs(3485)) or (layer2_outputs(7777));
    outputs(2926) <= layer2_outputs(3788);
    outputs(2927) <= not(layer2_outputs(7728));
    outputs(2928) <= not(layer2_outputs(2970)) or (layer2_outputs(6775));
    outputs(2929) <= not(layer2_outputs(5424));
    outputs(2930) <= layer2_outputs(4755);
    outputs(2931) <= layer2_outputs(6479);
    outputs(2932) <= not(layer2_outputs(6596));
    outputs(2933) <= not(layer2_outputs(7724));
    outputs(2934) <= (layer2_outputs(6279)) xor (layer2_outputs(5016));
    outputs(2935) <= not((layer2_outputs(1855)) xor (layer2_outputs(6267)));
    outputs(2936) <= layer2_outputs(8061);
    outputs(2937) <= (layer2_outputs(6646)) xor (layer2_outputs(1450));
    outputs(2938) <= layer2_outputs(5699);
    outputs(2939) <= layer2_outputs(9632);
    outputs(2940) <= not((layer2_outputs(7362)) and (layer2_outputs(4115)));
    outputs(2941) <= layer2_outputs(8854);
    outputs(2942) <= (layer2_outputs(4298)) xor (layer2_outputs(2683));
    outputs(2943) <= not(layer2_outputs(8453));
    outputs(2944) <= not(layer2_outputs(937));
    outputs(2945) <= not(layer2_outputs(299));
    outputs(2946) <= not(layer2_outputs(2260)) or (layer2_outputs(4540));
    outputs(2947) <= (layer2_outputs(2044)) xor (layer2_outputs(5864));
    outputs(2948) <= not(layer2_outputs(5713));
    outputs(2949) <= not(layer2_outputs(1504));
    outputs(2950) <= not((layer2_outputs(185)) or (layer2_outputs(3500)));
    outputs(2951) <= (layer2_outputs(3712)) xor (layer2_outputs(3294));
    outputs(2952) <= not((layer2_outputs(2495)) xor (layer2_outputs(3270)));
    outputs(2953) <= layer2_outputs(5082);
    outputs(2954) <= layer2_outputs(3789);
    outputs(2955) <= not(layer2_outputs(2205));
    outputs(2956) <= not(layer2_outputs(4078));
    outputs(2957) <= not(layer2_outputs(10008));
    outputs(2958) <= (layer2_outputs(8015)) and not (layer2_outputs(2138));
    outputs(2959) <= layer2_outputs(1207);
    outputs(2960) <= not(layer2_outputs(7518)) or (layer2_outputs(6251));
    outputs(2961) <= not(layer2_outputs(4708));
    outputs(2962) <= layer2_outputs(7939);
    outputs(2963) <= not(layer2_outputs(2241)) or (layer2_outputs(649));
    outputs(2964) <= (layer2_outputs(8254)) and (layer2_outputs(6308));
    outputs(2965) <= not((layer2_outputs(3702)) and (layer2_outputs(6783)));
    outputs(2966) <= not((layer2_outputs(8974)) xor (layer2_outputs(6657)));
    outputs(2967) <= layer2_outputs(2756);
    outputs(2968) <= not(layer2_outputs(3046));
    outputs(2969) <= not(layer2_outputs(6696));
    outputs(2970) <= (layer2_outputs(7357)) or (layer2_outputs(2259));
    outputs(2971) <= layer2_outputs(9275);
    outputs(2972) <= layer2_outputs(8906);
    outputs(2973) <= layer2_outputs(6790);
    outputs(2974) <= not(layer2_outputs(248));
    outputs(2975) <= not(layer2_outputs(2218));
    outputs(2976) <= not((layer2_outputs(5983)) xor (layer2_outputs(7412)));
    outputs(2977) <= not(layer2_outputs(8849));
    outputs(2978) <= (layer2_outputs(115)) and not (layer2_outputs(10233));
    outputs(2979) <= not(layer2_outputs(2222));
    outputs(2980) <= not(layer2_outputs(2211)) or (layer2_outputs(7106));
    outputs(2981) <= layer2_outputs(7926);
    outputs(2982) <= layer2_outputs(5626);
    outputs(2983) <= not(layer2_outputs(2270));
    outputs(2984) <= not(layer2_outputs(4049));
    outputs(2985) <= layer2_outputs(7605);
    outputs(2986) <= layer2_outputs(8753);
    outputs(2987) <= not(layer2_outputs(3277));
    outputs(2988) <= layer2_outputs(7705);
    outputs(2989) <= layer2_outputs(477);
    outputs(2990) <= (layer2_outputs(6754)) or (layer2_outputs(8756));
    outputs(2991) <= (layer2_outputs(1890)) xor (layer2_outputs(4921));
    outputs(2992) <= layer2_outputs(4557);
    outputs(2993) <= (layer2_outputs(4902)) xor (layer2_outputs(7987));
    outputs(2994) <= layer2_outputs(63);
    outputs(2995) <= not((layer2_outputs(3337)) xor (layer2_outputs(1999)));
    outputs(2996) <= layer2_outputs(7137);
    outputs(2997) <= not((layer2_outputs(5746)) or (layer2_outputs(929)));
    outputs(2998) <= not(layer2_outputs(8083)) or (layer2_outputs(3142));
    outputs(2999) <= not(layer2_outputs(428));
    outputs(3000) <= not(layer2_outputs(3500));
    outputs(3001) <= not(layer2_outputs(5370));
    outputs(3002) <= not(layer2_outputs(2910));
    outputs(3003) <= layer2_outputs(101);
    outputs(3004) <= not(layer2_outputs(9259));
    outputs(3005) <= layer2_outputs(6957);
    outputs(3006) <= not((layer2_outputs(9509)) xor (layer2_outputs(8608)));
    outputs(3007) <= not(layer2_outputs(5287));
    outputs(3008) <= (layer2_outputs(8728)) and not (layer2_outputs(6801));
    outputs(3009) <= (layer2_outputs(395)) and not (layer2_outputs(6858));
    outputs(3010) <= not(layer2_outputs(3147));
    outputs(3011) <= layer2_outputs(4028);
    outputs(3012) <= layer2_outputs(4160);
    outputs(3013) <= layer2_outputs(2705);
    outputs(3014) <= (layer2_outputs(77)) and not (layer2_outputs(4959));
    outputs(3015) <= not(layer2_outputs(4585));
    outputs(3016) <= not((layer2_outputs(550)) and (layer2_outputs(3926)));
    outputs(3017) <= not(layer2_outputs(5896));
    outputs(3018) <= (layer2_outputs(5921)) and not (layer2_outputs(9731));
    outputs(3019) <= (layer2_outputs(4588)) and not (layer2_outputs(3286));
    outputs(3020) <= not(layer2_outputs(4246)) or (layer2_outputs(563));
    outputs(3021) <= layer2_outputs(9616);
    outputs(3022) <= (layer2_outputs(2998)) and not (layer2_outputs(4906));
    outputs(3023) <= not(layer2_outputs(942)) or (layer2_outputs(1831));
    outputs(3024) <= not(layer2_outputs(349));
    outputs(3025) <= (layer2_outputs(394)) and not (layer2_outputs(3497));
    outputs(3026) <= not(layer2_outputs(1132));
    outputs(3027) <= (layer2_outputs(5917)) and not (layer2_outputs(96));
    outputs(3028) <= layer2_outputs(3696);
    outputs(3029) <= not(layer2_outputs(3007));
    outputs(3030) <= not(layer2_outputs(316)) or (layer2_outputs(368));
    outputs(3031) <= (layer2_outputs(998)) and (layer2_outputs(2996));
    outputs(3032) <= (layer2_outputs(7128)) or (layer2_outputs(2360));
    outputs(3033) <= not(layer2_outputs(2239));
    outputs(3034) <= not(layer2_outputs(4196));
    outputs(3035) <= not(layer2_outputs(5608));
    outputs(3036) <= layer2_outputs(464);
    outputs(3037) <= (layer2_outputs(9450)) and (layer2_outputs(7133));
    outputs(3038) <= layer2_outputs(2687);
    outputs(3039) <= layer2_outputs(1786);
    outputs(3040) <= not((layer2_outputs(136)) and (layer2_outputs(3584)));
    outputs(3041) <= (layer2_outputs(2377)) and (layer2_outputs(3023));
    outputs(3042) <= not(layer2_outputs(2435));
    outputs(3043) <= (layer2_outputs(6792)) or (layer2_outputs(1837));
    outputs(3044) <= layer2_outputs(4605);
    outputs(3045) <= not((layer2_outputs(2972)) or (layer2_outputs(7279)));
    outputs(3046) <= not((layer2_outputs(4273)) or (layer2_outputs(9714)));
    outputs(3047) <= not(layer2_outputs(8234));
    outputs(3048) <= not(layer2_outputs(2100)) or (layer2_outputs(5611));
    outputs(3049) <= not(layer2_outputs(6349));
    outputs(3050) <= not(layer2_outputs(9025));
    outputs(3051) <= layer2_outputs(4919);
    outputs(3052) <= (layer2_outputs(1224)) and (layer2_outputs(8251));
    outputs(3053) <= not(layer2_outputs(9986));
    outputs(3054) <= (layer2_outputs(632)) and not (layer2_outputs(6698));
    outputs(3055) <= not(layer2_outputs(2557));
    outputs(3056) <= not(layer2_outputs(5518));
    outputs(3057) <= (layer2_outputs(4191)) and (layer2_outputs(9122));
    outputs(3058) <= not((layer2_outputs(4016)) xor (layer2_outputs(5294)));
    outputs(3059) <= layer2_outputs(6204);
    outputs(3060) <= (layer2_outputs(7167)) xor (layer2_outputs(4834));
    outputs(3061) <= not(layer2_outputs(3880)) or (layer2_outputs(10073));
    outputs(3062) <= not((layer2_outputs(4562)) and (layer2_outputs(994)));
    outputs(3063) <= not(layer2_outputs(6278));
    outputs(3064) <= layer2_outputs(502);
    outputs(3065) <= not(layer2_outputs(4420)) or (layer2_outputs(9197));
    outputs(3066) <= layer2_outputs(9821);
    outputs(3067) <= not(layer2_outputs(8232));
    outputs(3068) <= not(layer2_outputs(8075));
    outputs(3069) <= layer2_outputs(6461);
    outputs(3070) <= layer2_outputs(7993);
    outputs(3071) <= layer2_outputs(2641);
    outputs(3072) <= not(layer2_outputs(3799));
    outputs(3073) <= layer2_outputs(7277);
    outputs(3074) <= not((layer2_outputs(7255)) xor (layer2_outputs(873)));
    outputs(3075) <= not(layer2_outputs(2332));
    outputs(3076) <= layer2_outputs(7392);
    outputs(3077) <= not((layer2_outputs(1362)) xor (layer2_outputs(7727)));
    outputs(3078) <= layer2_outputs(7278);
    outputs(3079) <= not((layer2_outputs(2370)) xor (layer2_outputs(5049)));
    outputs(3080) <= (layer2_outputs(5956)) and (layer2_outputs(385));
    outputs(3081) <= not((layer2_outputs(9089)) or (layer2_outputs(9179)));
    outputs(3082) <= layer2_outputs(6400);
    outputs(3083) <= not(layer2_outputs(8355));
    outputs(3084) <= not(layer2_outputs(5341));
    outputs(3085) <= layer2_outputs(3430);
    outputs(3086) <= layer2_outputs(3068);
    outputs(3087) <= not(layer2_outputs(5899));
    outputs(3088) <= (layer2_outputs(6501)) and not (layer2_outputs(7486));
    outputs(3089) <= (layer2_outputs(9247)) and not (layer2_outputs(2873));
    outputs(3090) <= layer2_outputs(2577);
    outputs(3091) <= not(layer2_outputs(1394));
    outputs(3092) <= (layer2_outputs(482)) and (layer2_outputs(6281));
    outputs(3093) <= layer2_outputs(3850);
    outputs(3094) <= layer2_outputs(3940);
    outputs(3095) <= not(layer2_outputs(7697));
    outputs(3096) <= (layer2_outputs(1764)) and not (layer2_outputs(3678));
    outputs(3097) <= not((layer2_outputs(5413)) xor (layer2_outputs(2748)));
    outputs(3098) <= layer2_outputs(148);
    outputs(3099) <= not(layer2_outputs(4016));
    outputs(3100) <= (layer2_outputs(1599)) and not (layer2_outputs(7733));
    outputs(3101) <= (layer2_outputs(5253)) and (layer2_outputs(1442));
    outputs(3102) <= layer2_outputs(8915);
    outputs(3103) <= layer2_outputs(2449);
    outputs(3104) <= layer2_outputs(3494);
    outputs(3105) <= not(layer2_outputs(4498)) or (layer2_outputs(5344));
    outputs(3106) <= not(layer2_outputs(1550));
    outputs(3107) <= not(layer2_outputs(3847));
    outputs(3108) <= not(layer2_outputs(7527));
    outputs(3109) <= layer2_outputs(9071);
    outputs(3110) <= not(layer2_outputs(3336));
    outputs(3111) <= layer2_outputs(9517);
    outputs(3112) <= not(layer2_outputs(663));
    outputs(3113) <= not(layer2_outputs(9098));
    outputs(3114) <= layer2_outputs(8390);
    outputs(3115) <= layer2_outputs(5061);
    outputs(3116) <= layer2_outputs(5025);
    outputs(3117) <= not(layer2_outputs(8716)) or (layer2_outputs(8231));
    outputs(3118) <= layer2_outputs(1781);
    outputs(3119) <= layer2_outputs(1974);
    outputs(3120) <= layer2_outputs(320);
    outputs(3121) <= not(layer2_outputs(9550));
    outputs(3122) <= (layer2_outputs(1423)) xor (layer2_outputs(4242));
    outputs(3123) <= (layer2_outputs(7139)) and (layer2_outputs(1104));
    outputs(3124) <= not((layer2_outputs(3205)) xor (layer2_outputs(7409)));
    outputs(3125) <= not(layer2_outputs(1850));
    outputs(3126) <= (layer2_outputs(9999)) xor (layer2_outputs(4106));
    outputs(3127) <= layer2_outputs(8012);
    outputs(3128) <= not(layer2_outputs(9872));
    outputs(3129) <= not(layer2_outputs(3544));
    outputs(3130) <= layer2_outputs(3202);
    outputs(3131) <= layer2_outputs(7847);
    outputs(3132) <= not(layer2_outputs(8908)) or (layer2_outputs(1121));
    outputs(3133) <= (layer2_outputs(6297)) xor (layer2_outputs(9771));
    outputs(3134) <= not(layer2_outputs(2688)) or (layer2_outputs(1343));
    outputs(3135) <= not(layer2_outputs(10214)) or (layer2_outputs(10166));
    outputs(3136) <= not(layer2_outputs(2223));
    outputs(3137) <= not(layer2_outputs(7384));
    outputs(3138) <= (layer2_outputs(9887)) xor (layer2_outputs(3314));
    outputs(3139) <= layer2_outputs(364);
    outputs(3140) <= layer2_outputs(8128);
    outputs(3141) <= not(layer2_outputs(9555));
    outputs(3142) <= layer2_outputs(3413);
    outputs(3143) <= not((layer2_outputs(6374)) or (layer2_outputs(3909)));
    outputs(3144) <= not(layer2_outputs(6625));
    outputs(3145) <= layer2_outputs(1577);
    outputs(3146) <= layer2_outputs(4609);
    outputs(3147) <= not(layer2_outputs(1118));
    outputs(3148) <= (layer2_outputs(4482)) and not (layer2_outputs(9716));
    outputs(3149) <= not(layer2_outputs(5830)) or (layer2_outputs(9580));
    outputs(3150) <= not(layer2_outputs(9572));
    outputs(3151) <= not((layer2_outputs(8394)) xor (layer2_outputs(7067)));
    outputs(3152) <= not(layer2_outputs(1836));
    outputs(3153) <= not(layer2_outputs(6242));
    outputs(3154) <= not(layer2_outputs(2019)) or (layer2_outputs(7910));
    outputs(3155) <= layer2_outputs(7886);
    outputs(3156) <= (layer2_outputs(4010)) or (layer2_outputs(8224));
    outputs(3157) <= not((layer2_outputs(1866)) xor (layer2_outputs(8299)));
    outputs(3158) <= (layer2_outputs(8747)) and (layer2_outputs(8797));
    outputs(3159) <= layer2_outputs(1588);
    outputs(3160) <= not(layer2_outputs(2656));
    outputs(3161) <= not(layer2_outputs(8613));
    outputs(3162) <= not(layer2_outputs(6477));
    outputs(3163) <= not(layer2_outputs(2987));
    outputs(3164) <= not(layer2_outputs(2274));
    outputs(3165) <= layer2_outputs(8397);
    outputs(3166) <= not(layer2_outputs(5395));
    outputs(3167) <= layer2_outputs(5829);
    outputs(3168) <= layer2_outputs(1827);
    outputs(3169) <= (layer2_outputs(5381)) and (layer2_outputs(4739));
    outputs(3170) <= (layer2_outputs(2191)) and not (layer2_outputs(8735));
    outputs(3171) <= not(layer2_outputs(6601));
    outputs(3172) <= not(layer2_outputs(1890));
    outputs(3173) <= (layer2_outputs(2651)) and not (layer2_outputs(3061));
    outputs(3174) <= (layer2_outputs(1247)) and (layer2_outputs(2561));
    outputs(3175) <= not(layer2_outputs(6135));
    outputs(3176) <= (layer2_outputs(9420)) xor (layer2_outputs(9049));
    outputs(3177) <= not((layer2_outputs(187)) xor (layer2_outputs(9662)));
    outputs(3178) <= layer2_outputs(158);
    outputs(3179) <= (layer2_outputs(9668)) and not (layer2_outputs(10075));
    outputs(3180) <= layer2_outputs(4754);
    outputs(3181) <= layer2_outputs(9484);
    outputs(3182) <= not(layer2_outputs(7608));
    outputs(3183) <= (layer2_outputs(321)) and not (layer2_outputs(2127));
    outputs(3184) <= not((layer2_outputs(9283)) xor (layer2_outputs(8310)));
    outputs(3185) <= (layer2_outputs(6820)) xor (layer2_outputs(6989));
    outputs(3186) <= (layer2_outputs(3468)) and (layer2_outputs(7688));
    outputs(3187) <= layer2_outputs(6730);
    outputs(3188) <= not(layer2_outputs(4279));
    outputs(3189) <= not(layer2_outputs(3962));
    outputs(3190) <= (layer2_outputs(4307)) and not (layer2_outputs(872));
    outputs(3191) <= layer2_outputs(6567);
    outputs(3192) <= (layer2_outputs(9814)) and (layer2_outputs(5385));
    outputs(3193) <= not(layer2_outputs(9040)) or (layer2_outputs(4887));
    outputs(3194) <= layer2_outputs(3018);
    outputs(3195) <= not(layer2_outputs(4499));
    outputs(3196) <= not(layer2_outputs(6933));
    outputs(3197) <= not(layer2_outputs(5262));
    outputs(3198) <= layer2_outputs(4263);
    outputs(3199) <= not((layer2_outputs(4390)) xor (layer2_outputs(2277)));
    outputs(3200) <= (layer2_outputs(2883)) xor (layer2_outputs(2916));
    outputs(3201) <= (layer2_outputs(7589)) xor (layer2_outputs(3380));
    outputs(3202) <= not(layer2_outputs(2986));
    outputs(3203) <= (layer2_outputs(7122)) and (layer2_outputs(500));
    outputs(3204) <= not(layer2_outputs(4271));
    outputs(3205) <= not((layer2_outputs(5340)) and (layer2_outputs(8335)));
    outputs(3206) <= not(layer2_outputs(1565));
    outputs(3207) <= not(layer2_outputs(1788));
    outputs(3208) <= layer2_outputs(7969);
    outputs(3209) <= layer2_outputs(1190);
    outputs(3210) <= not(layer2_outputs(3084));
    outputs(3211) <= not(layer2_outputs(7686));
    outputs(3212) <= (layer2_outputs(1)) or (layer2_outputs(9638));
    outputs(3213) <= (layer2_outputs(9257)) xor (layer2_outputs(896));
    outputs(3214) <= (layer2_outputs(2487)) and not (layer2_outputs(1449));
    outputs(3215) <= not(layer2_outputs(9826));
    outputs(3216) <= layer2_outputs(6902);
    outputs(3217) <= layer2_outputs(4725);
    outputs(3218) <= not(layer2_outputs(2999));
    outputs(3219) <= (layer2_outputs(912)) or (layer2_outputs(2851));
    outputs(3220) <= not((layer2_outputs(3491)) xor (layer2_outputs(5714)));
    outputs(3221) <= (layer2_outputs(1961)) and (layer2_outputs(8688));
    outputs(3222) <= not((layer2_outputs(4917)) xor (layer2_outputs(4103)));
    outputs(3223) <= not((layer2_outputs(5562)) xor (layer2_outputs(308)));
    outputs(3224) <= not((layer2_outputs(2977)) xor (layer2_outputs(7389)));
    outputs(3225) <= layer2_outputs(604);
    outputs(3226) <= not((layer2_outputs(7243)) xor (layer2_outputs(4973)));
    outputs(3227) <= layer2_outputs(5827);
    outputs(3228) <= layer2_outputs(9537);
    outputs(3229) <= not((layer2_outputs(9915)) xor (layer2_outputs(2980)));
    outputs(3230) <= not((layer2_outputs(5511)) or (layer2_outputs(7367)));
    outputs(3231) <= not((layer2_outputs(4405)) xor (layer2_outputs(2211)));
    outputs(3232) <= (layer2_outputs(1222)) xor (layer2_outputs(5779));
    outputs(3233) <= not((layer2_outputs(3528)) or (layer2_outputs(5957)));
    outputs(3234) <= not(layer2_outputs(6594));
    outputs(3235) <= not((layer2_outputs(6532)) xor (layer2_outputs(393)));
    outputs(3236) <= not((layer2_outputs(1657)) and (layer2_outputs(9928)));
    outputs(3237) <= layer2_outputs(8521);
    outputs(3238) <= not((layer2_outputs(8385)) xor (layer2_outputs(1448)));
    outputs(3239) <= (layer2_outputs(7360)) and not (layer2_outputs(9987));
    outputs(3240) <= layer2_outputs(7888);
    outputs(3241) <= not((layer2_outputs(7431)) xor (layer2_outputs(730)));
    outputs(3242) <= layer2_outputs(1802);
    outputs(3243) <= not(layer2_outputs(10174)) or (layer2_outputs(1463));
    outputs(3244) <= layer2_outputs(7392);
    outputs(3245) <= (layer2_outputs(4679)) xor (layer2_outputs(6057));
    outputs(3246) <= (layer2_outputs(4458)) and not (layer2_outputs(7902));
    outputs(3247) <= layer2_outputs(4291);
    outputs(3248) <= (layer2_outputs(4165)) and (layer2_outputs(8254));
    outputs(3249) <= not(layer2_outputs(4518));
    outputs(3250) <= not((layer2_outputs(3661)) xor (layer2_outputs(8117)));
    outputs(3251) <= not((layer2_outputs(9594)) xor (layer2_outputs(6855)));
    outputs(3252) <= (layer2_outputs(3047)) and not (layer2_outputs(3530));
    outputs(3253) <= (layer2_outputs(9893)) or (layer2_outputs(742));
    outputs(3254) <= not(layer2_outputs(6175));
    outputs(3255) <= layer2_outputs(8255);
    outputs(3256) <= (layer2_outputs(9897)) xor (layer2_outputs(9387));
    outputs(3257) <= layer2_outputs(7704);
    outputs(3258) <= (layer2_outputs(5974)) and not (layer2_outputs(4678));
    outputs(3259) <= (layer2_outputs(5767)) xor (layer2_outputs(8465));
    outputs(3260) <= not((layer2_outputs(6877)) xor (layer2_outputs(9445)));
    outputs(3261) <= not((layer2_outputs(5215)) xor (layer2_outputs(8717)));
    outputs(3262) <= layer2_outputs(5948);
    outputs(3263) <= not(layer2_outputs(984)) or (layer2_outputs(1864));
    outputs(3264) <= not((layer2_outputs(4634)) and (layer2_outputs(8901)));
    outputs(3265) <= not(layer2_outputs(6465));
    outputs(3266) <= layer2_outputs(4541);
    outputs(3267) <= not(layer2_outputs(4552));
    outputs(3268) <= layer2_outputs(6430);
    outputs(3269) <= (layer2_outputs(3141)) and not (layer2_outputs(190));
    outputs(3270) <= not(layer2_outputs(40));
    outputs(3271) <= not(layer2_outputs(2202));
    outputs(3272) <= (layer2_outputs(9412)) and (layer2_outputs(6478));
    outputs(3273) <= layer2_outputs(2490);
    outputs(3274) <= (layer2_outputs(3575)) xor (layer2_outputs(9920));
    outputs(3275) <= layer2_outputs(4997);
    outputs(3276) <= not(layer2_outputs(9432));
    outputs(3277) <= not(layer2_outputs(1443)) or (layer2_outputs(9160));
    outputs(3278) <= not((layer2_outputs(4473)) xor (layer2_outputs(6918)));
    outputs(3279) <= not(layer2_outputs(728)) or (layer2_outputs(7729));
    outputs(3280) <= not((layer2_outputs(1368)) xor (layer2_outputs(3922)));
    outputs(3281) <= layer2_outputs(10144);
    outputs(3282) <= not(layer2_outputs(3634));
    outputs(3283) <= layer2_outputs(2851);
    outputs(3284) <= (layer2_outputs(480)) and not (layer2_outputs(2970));
    outputs(3285) <= not(layer2_outputs(8496));
    outputs(3286) <= layer2_outputs(5460);
    outputs(3287) <= not(layer2_outputs(6583)) or (layer2_outputs(5692));
    outputs(3288) <= (layer2_outputs(2909)) xor (layer2_outputs(287));
    outputs(3289) <= not(layer2_outputs(9300));
    outputs(3290) <= layer2_outputs(2838);
    outputs(3291) <= layer2_outputs(3621);
    outputs(3292) <= layer2_outputs(10208);
    outputs(3293) <= not((layer2_outputs(3861)) xor (layer2_outputs(7426)));
    outputs(3294) <= not(layer2_outputs(4112));
    outputs(3295) <= not((layer2_outputs(4444)) xor (layer2_outputs(3134)));
    outputs(3296) <= not(layer2_outputs(280));
    outputs(3297) <= not((layer2_outputs(6456)) xor (layer2_outputs(2122)));
    outputs(3298) <= layer2_outputs(5720);
    outputs(3299) <= (layer2_outputs(5752)) xor (layer2_outputs(6762));
    outputs(3300) <= layer2_outputs(6603);
    outputs(3301) <= not((layer2_outputs(7221)) xor (layer2_outputs(8325)));
    outputs(3302) <= not((layer2_outputs(6921)) or (layer2_outputs(9769)));
    outputs(3303) <= not((layer2_outputs(7996)) xor (layer2_outputs(7460)));
    outputs(3304) <= (layer2_outputs(3960)) xor (layer2_outputs(876));
    outputs(3305) <= (layer2_outputs(7859)) and not (layer2_outputs(8615));
    outputs(3306) <= (layer2_outputs(282)) xor (layer2_outputs(5920));
    outputs(3307) <= not(layer2_outputs(5968));
    outputs(3308) <= not((layer2_outputs(3473)) or (layer2_outputs(1748)));
    outputs(3309) <= (layer2_outputs(8004)) xor (layer2_outputs(2928));
    outputs(3310) <= not(layer2_outputs(8061)) or (layer2_outputs(9725));
    outputs(3311) <= not(layer2_outputs(2551));
    outputs(3312) <= (layer2_outputs(5076)) xor (layer2_outputs(8217));
    outputs(3313) <= not((layer2_outputs(2815)) xor (layer2_outputs(1935)));
    outputs(3314) <= not(layer2_outputs(54));
    outputs(3315) <= (layer2_outputs(4063)) and not (layer2_outputs(4395));
    outputs(3316) <= layer2_outputs(5502);
    outputs(3317) <= not(layer2_outputs(9094));
    outputs(3318) <= not((layer2_outputs(3728)) xor (layer2_outputs(10063)));
    outputs(3319) <= not(layer2_outputs(294));
    outputs(3320) <= not(layer2_outputs(6629));
    outputs(3321) <= layer2_outputs(8158);
    outputs(3322) <= not((layer2_outputs(6319)) and (layer2_outputs(8529)));
    outputs(3323) <= not(layer2_outputs(2333)) or (layer2_outputs(1501));
    outputs(3324) <= (layer2_outputs(4144)) xor (layer2_outputs(8798));
    outputs(3325) <= (layer2_outputs(6162)) xor (layer2_outputs(964));
    outputs(3326) <= not(layer2_outputs(1772));
    outputs(3327) <= not(layer2_outputs(6343));
    outputs(3328) <= not(layer2_outputs(6613));
    outputs(3329) <= (layer2_outputs(5322)) xor (layer2_outputs(9385));
    outputs(3330) <= (layer2_outputs(2792)) and not (layer2_outputs(3098));
    outputs(3331) <= layer2_outputs(4323);
    outputs(3332) <= not(layer2_outputs(617)) or (layer2_outputs(2095));
    outputs(3333) <= not(layer2_outputs(3076));
    outputs(3334) <= layer2_outputs(3052);
    outputs(3335) <= (layer2_outputs(9634)) xor (layer2_outputs(5272));
    outputs(3336) <= not(layer2_outputs(811));
    outputs(3337) <= layer2_outputs(3211);
    outputs(3338) <= layer2_outputs(706);
    outputs(3339) <= (layer2_outputs(9200)) xor (layer2_outputs(9083));
    outputs(3340) <= not(layer2_outputs(9734));
    outputs(3341) <= layer2_outputs(8826);
    outputs(3342) <= not(layer2_outputs(8603));
    outputs(3343) <= (layer2_outputs(3935)) and (layer2_outputs(4621));
    outputs(3344) <= layer2_outputs(9921);
    outputs(3345) <= layer2_outputs(4936);
    outputs(3346) <= layer2_outputs(9115);
    outputs(3347) <= (layer2_outputs(4809)) and not (layer2_outputs(8919));
    outputs(3348) <= (layer2_outputs(4672)) xor (layer2_outputs(4592));
    outputs(3349) <= (layer2_outputs(3492)) xor (layer2_outputs(7832));
    outputs(3350) <= not(layer2_outputs(9462));
    outputs(3351) <= layer2_outputs(7820);
    outputs(3352) <= (layer2_outputs(9197)) and not (layer2_outputs(5945));
    outputs(3353) <= not(layer2_outputs(8603));
    outputs(3354) <= layer2_outputs(2584);
    outputs(3355) <= (layer2_outputs(4402)) xor (layer2_outputs(8060));
    outputs(3356) <= not((layer2_outputs(4169)) xor (layer2_outputs(2931)));
    outputs(3357) <= (layer2_outputs(1163)) xor (layer2_outputs(3186));
    outputs(3358) <= not(layer2_outputs(2013));
    outputs(3359) <= not(layer2_outputs(1962));
    outputs(3360) <= layer2_outputs(10005);
    outputs(3361) <= (layer2_outputs(4388)) xor (layer2_outputs(2201));
    outputs(3362) <= layer2_outputs(4804);
    outputs(3363) <= not((layer2_outputs(9206)) xor (layer2_outputs(8063)));
    outputs(3364) <= not(layer2_outputs(5878));
    outputs(3365) <= (layer2_outputs(6607)) and not (layer2_outputs(346));
    outputs(3366) <= (layer2_outputs(1807)) and not (layer2_outputs(6168));
    outputs(3367) <= not(layer2_outputs(6349));
    outputs(3368) <= not(layer2_outputs(7524));
    outputs(3369) <= layer2_outputs(8985);
    outputs(3370) <= not(layer2_outputs(5263)) or (layer2_outputs(985));
    outputs(3371) <= (layer2_outputs(4796)) xor (layer2_outputs(6728));
    outputs(3372) <= (layer2_outputs(1902)) xor (layer2_outputs(1440));
    outputs(3373) <= not((layer2_outputs(8808)) xor (layer2_outputs(7311)));
    outputs(3374) <= layer2_outputs(1758);
    outputs(3375) <= not(layer2_outputs(7452));
    outputs(3376) <= layer2_outputs(5545);
    outputs(3377) <= not((layer2_outputs(9219)) or (layer2_outputs(4485)));
    outputs(3378) <= not(layer2_outputs(8306)) or (layer2_outputs(9719));
    outputs(3379) <= not(layer2_outputs(1565));
    outputs(3380) <= layer2_outputs(540);
    outputs(3381) <= (layer2_outputs(911)) and (layer2_outputs(5043));
    outputs(3382) <= not(layer2_outputs(3842));
    outputs(3383) <= (layer2_outputs(10079)) or (layer2_outputs(1017));
    outputs(3384) <= layer2_outputs(7847);
    outputs(3385) <= not(layer2_outputs(1808));
    outputs(3386) <= not((layer2_outputs(5353)) xor (layer2_outputs(9996)));
    outputs(3387) <= not(layer2_outputs(3006));
    outputs(3388) <= not((layer2_outputs(5664)) xor (layer2_outputs(6376)));
    outputs(3389) <= (layer2_outputs(9063)) and (layer2_outputs(10232));
    outputs(3390) <= (layer2_outputs(1270)) xor (layer2_outputs(6150));
    outputs(3391) <= layer2_outputs(3426);
    outputs(3392) <= not((layer2_outputs(9727)) xor (layer2_outputs(4890)));
    outputs(3393) <= not(layer2_outputs(8009));
    outputs(3394) <= not(layer2_outputs(1814));
    outputs(3395) <= not(layer2_outputs(1217));
    outputs(3396) <= not((layer2_outputs(6443)) xor (layer2_outputs(4333)));
    outputs(3397) <= not(layer2_outputs(3345));
    outputs(3398) <= layer2_outputs(7905);
    outputs(3399) <= (layer2_outputs(10130)) and not (layer2_outputs(836));
    outputs(3400) <= (layer2_outputs(1554)) and not (layer2_outputs(5759));
    outputs(3401) <= layer2_outputs(7738);
    outputs(3402) <= not(layer2_outputs(5719));
    outputs(3403) <= layer2_outputs(3981);
    outputs(3404) <= not(layer2_outputs(4103));
    outputs(3405) <= not((layer2_outputs(9225)) xor (layer2_outputs(643)));
    outputs(3406) <= (layer2_outputs(3372)) xor (layer2_outputs(870));
    outputs(3407) <= layer2_outputs(171);
    outputs(3408) <= layer2_outputs(1571);
    outputs(3409) <= layer2_outputs(7927);
    outputs(3410) <= not(layer2_outputs(3860));
    outputs(3411) <= not(layer2_outputs(2094));
    outputs(3412) <= (layer2_outputs(1075)) and not (layer2_outputs(8549));
    outputs(3413) <= (layer2_outputs(8602)) xor (layer2_outputs(7880));
    outputs(3414) <= layer2_outputs(10207);
    outputs(3415) <= layer2_outputs(9898);
    outputs(3416) <= not(layer2_outputs(6090));
    outputs(3417) <= not(layer2_outputs(6096)) or (layer2_outputs(7163));
    outputs(3418) <= not(layer2_outputs(354));
    outputs(3419) <= not((layer2_outputs(7707)) xor (layer2_outputs(7005)));
    outputs(3420) <= not((layer2_outputs(1642)) xor (layer2_outputs(3036)));
    outputs(3421) <= not(layer2_outputs(2140)) or (layer2_outputs(5625));
    outputs(3422) <= (layer2_outputs(7416)) and not (layer2_outputs(6309));
    outputs(3423) <= (layer2_outputs(9426)) or (layer2_outputs(5826));
    outputs(3424) <= not((layer2_outputs(8956)) xor (layer2_outputs(4387)));
    outputs(3425) <= not(layer2_outputs(4314));
    outputs(3426) <= not((layer2_outputs(1899)) xor (layer2_outputs(1912)));
    outputs(3427) <= not(layer2_outputs(23));
    outputs(3428) <= layer2_outputs(5110);
    outputs(3429) <= (layer2_outputs(7909)) and not (layer2_outputs(2364));
    outputs(3430) <= not(layer2_outputs(8124));
    outputs(3431) <= not(layer2_outputs(3343)) or (layer2_outputs(199));
    outputs(3432) <= not(layer2_outputs(9440));
    outputs(3433) <= (layer2_outputs(449)) and (layer2_outputs(5953));
    outputs(3434) <= layer2_outputs(5288);
    outputs(3435) <= not(layer2_outputs(286));
    outputs(3436) <= (layer2_outputs(6981)) and (layer2_outputs(8669));
    outputs(3437) <= not(layer2_outputs(1105));
    outputs(3438) <= not(layer2_outputs(5137));
    outputs(3439) <= layer2_outputs(5876);
    outputs(3440) <= not(layer2_outputs(5981));
    outputs(3441) <= layer2_outputs(3338);
    outputs(3442) <= layer2_outputs(988);
    outputs(3443) <= not(layer2_outputs(8475));
    outputs(3444) <= not((layer2_outputs(5391)) xor (layer2_outputs(5022)));
    outputs(3445) <= not(layer2_outputs(4992));
    outputs(3446) <= (layer2_outputs(9315)) and not (layer2_outputs(8770));
    outputs(3447) <= not(layer2_outputs(5546));
    outputs(3448) <= not(layer2_outputs(6961));
    outputs(3449) <= not(layer2_outputs(938));
    outputs(3450) <= layer2_outputs(3047);
    outputs(3451) <= (layer2_outputs(1881)) xor (layer2_outputs(7359));
    outputs(3452) <= layer2_outputs(5232);
    outputs(3453) <= layer2_outputs(4893);
    outputs(3454) <= layer2_outputs(6482);
    outputs(3455) <= layer2_outputs(758);
    outputs(3456) <= not(layer2_outputs(9671));
    outputs(3457) <= not(layer2_outputs(8846));
    outputs(3458) <= layer2_outputs(8997);
    outputs(3459) <= (layer2_outputs(5279)) xor (layer2_outputs(7427));
    outputs(3460) <= layer2_outputs(8274);
    outputs(3461) <= (layer2_outputs(2917)) or (layer2_outputs(486));
    outputs(3462) <= (layer2_outputs(6214)) xor (layer2_outputs(8089));
    outputs(3463) <= not((layer2_outputs(8165)) xor (layer2_outputs(5791)));
    outputs(3464) <= (layer2_outputs(6691)) or (layer2_outputs(9322));
    outputs(3465) <= layer2_outputs(3870);
    outputs(3466) <= layer2_outputs(8952);
    outputs(3467) <= not((layer2_outputs(2531)) xor (layer2_outputs(4341)));
    outputs(3468) <= (layer2_outputs(4559)) xor (layer2_outputs(7541));
    outputs(3469) <= not((layer2_outputs(3037)) xor (layer2_outputs(2830)));
    outputs(3470) <= (layer2_outputs(3926)) and (layer2_outputs(3822));
    outputs(3471) <= (layer2_outputs(7278)) and not (layer2_outputs(8107));
    outputs(3472) <= not(layer2_outputs(9791));
    outputs(3473) <= layer2_outputs(10129);
    outputs(3474) <= (layer2_outputs(2158)) xor (layer2_outputs(4047));
    outputs(3475) <= not(layer2_outputs(7576));
    outputs(3476) <= layer2_outputs(8793);
    outputs(3477) <= layer2_outputs(337);
    outputs(3478) <= not(layer2_outputs(8177));
    outputs(3479) <= layer2_outputs(5835);
    outputs(3480) <= not(layer2_outputs(9516));
    outputs(3481) <= layer2_outputs(5775);
    outputs(3482) <= not(layer2_outputs(246)) or (layer2_outputs(2156));
    outputs(3483) <= not((layer2_outputs(7679)) xor (layer2_outputs(6145)));
    outputs(3484) <= (layer2_outputs(6832)) xor (layer2_outputs(10112));
    outputs(3485) <= (layer2_outputs(298)) and (layer2_outputs(4439));
    outputs(3486) <= (layer2_outputs(37)) or (layer2_outputs(1995));
    outputs(3487) <= not(layer2_outputs(4416)) or (layer2_outputs(3392));
    outputs(3488) <= not(layer2_outputs(901));
    outputs(3489) <= layer2_outputs(3952);
    outputs(3490) <= layer2_outputs(4541);
    outputs(3491) <= layer2_outputs(2801);
    outputs(3492) <= not((layer2_outputs(10027)) or (layer2_outputs(7015)));
    outputs(3493) <= layer2_outputs(3839);
    outputs(3494) <= layer2_outputs(877);
    outputs(3495) <= (layer2_outputs(2)) and not (layer2_outputs(2693));
    outputs(3496) <= (layer2_outputs(3899)) and (layer2_outputs(9536));
    outputs(3497) <= not((layer2_outputs(2981)) and (layer2_outputs(7033)));
    outputs(3498) <= not(layer2_outputs(10029));
    outputs(3499) <= not(layer2_outputs(4113));
    outputs(3500) <= layer2_outputs(8195);
    outputs(3501) <= (layer2_outputs(4140)) and (layer2_outputs(2262));
    outputs(3502) <= (layer2_outputs(2357)) or (layer2_outputs(5462));
    outputs(3503) <= not(layer2_outputs(2115));
    outputs(3504) <= (layer2_outputs(4665)) xor (layer2_outputs(3024));
    outputs(3505) <= (layer2_outputs(544)) and (layer2_outputs(3746));
    outputs(3506) <= not((layer2_outputs(2040)) xor (layer2_outputs(425)));
    outputs(3507) <= not(layer2_outputs(7249)) or (layer2_outputs(4410));
    outputs(3508) <= (layer2_outputs(9277)) and not (layer2_outputs(4090));
    outputs(3509) <= not(layer2_outputs(4669)) or (layer2_outputs(5575));
    outputs(3510) <= layer2_outputs(605);
    outputs(3511) <= not((layer2_outputs(8903)) xor (layer2_outputs(8849)));
    outputs(3512) <= not((layer2_outputs(7979)) xor (layer2_outputs(6860)));
    outputs(3513) <= not((layer2_outputs(5993)) xor (layer2_outputs(4999)));
    outputs(3514) <= not(layer2_outputs(5492));
    outputs(3515) <= layer2_outputs(9234);
    outputs(3516) <= not(layer2_outputs(8031));
    outputs(3517) <= not((layer2_outputs(8973)) xor (layer2_outputs(4221)));
    outputs(3518) <= not(layer2_outputs(8564)) or (layer2_outputs(3222));
    outputs(3519) <= (layer2_outputs(8483)) xor (layer2_outputs(5024));
    outputs(3520) <= not((layer2_outputs(3538)) xor (layer2_outputs(3608)));
    outputs(3521) <= not((layer2_outputs(1596)) xor (layer2_outputs(2927)));
    outputs(3522) <= layer2_outputs(586);
    outputs(3523) <= not((layer2_outputs(3130)) xor (layer2_outputs(2662)));
    outputs(3524) <= not(layer2_outputs(7086));
    outputs(3525) <= not(layer2_outputs(275));
    outputs(3526) <= layer2_outputs(7552);
    outputs(3527) <= not(layer2_outputs(636));
    outputs(3528) <= (layer2_outputs(7160)) xor (layer2_outputs(7668));
    outputs(3529) <= layer2_outputs(5613);
    outputs(3530) <= layer2_outputs(2728);
    outputs(3531) <= layer2_outputs(1744);
    outputs(3532) <= layer2_outputs(2628);
    outputs(3533) <= not((layer2_outputs(2597)) or (layer2_outputs(1651)));
    outputs(3534) <= not((layer2_outputs(4954)) xor (layer2_outputs(9581)));
    outputs(3535) <= (layer2_outputs(4977)) and not (layer2_outputs(4735));
    outputs(3536) <= (layer2_outputs(9334)) and (layer2_outputs(6385));
    outputs(3537) <= (layer2_outputs(8913)) and (layer2_outputs(6658));
    outputs(3538) <= (layer2_outputs(8688)) and not (layer2_outputs(869));
    outputs(3539) <= not(layer2_outputs(1321));
    outputs(3540) <= not(layer2_outputs(8319));
    outputs(3541) <= layer2_outputs(8833);
    outputs(3542) <= not(layer2_outputs(1408));
    outputs(3543) <= (layer2_outputs(2067)) and (layer2_outputs(6293));
    outputs(3544) <= not(layer2_outputs(4810));
    outputs(3545) <= not(layer2_outputs(3189)) or (layer2_outputs(559));
    outputs(3546) <= not(layer2_outputs(1130));
    outputs(3547) <= layer2_outputs(7267);
    outputs(3548) <= not(layer2_outputs(1606));
    outputs(3549) <= not(layer2_outputs(9443));
    outputs(3550) <= not(layer2_outputs(1883));
    outputs(3551) <= not((layer2_outputs(1762)) xor (layer2_outputs(4140)));
    outputs(3552) <= not(layer2_outputs(3239));
    outputs(3553) <= not(layer2_outputs(841)) or (layer2_outputs(2822));
    outputs(3554) <= not(layer2_outputs(9227));
    outputs(3555) <= (layer2_outputs(9071)) and (layer2_outputs(145));
    outputs(3556) <= (layer2_outputs(4046)) and not (layer2_outputs(1116));
    outputs(3557) <= not(layer2_outputs(1059));
    outputs(3558) <= not(layer2_outputs(7930)) or (layer2_outputs(6900));
    outputs(3559) <= (layer2_outputs(714)) and (layer2_outputs(4543));
    outputs(3560) <= not(layer2_outputs(6211));
    outputs(3561) <= (layer2_outputs(6040)) xor (layer2_outputs(5867));
    outputs(3562) <= not(layer2_outputs(30)) or (layer2_outputs(7901));
    outputs(3563) <= not(layer2_outputs(9454));
    outputs(3564) <= not((layer2_outputs(1473)) xor (layer2_outputs(1873)));
    outputs(3565) <= not((layer2_outputs(9468)) or (layer2_outputs(406)));
    outputs(3566) <= layer2_outputs(2960);
    outputs(3567) <= layer2_outputs(9721);
    outputs(3568) <= (layer2_outputs(178)) xor (layer2_outputs(8070));
    outputs(3569) <= (layer2_outputs(2229)) xor (layer2_outputs(1406));
    outputs(3570) <= layer2_outputs(1690);
    outputs(3571) <= (layer2_outputs(7174)) and not (layer2_outputs(4236));
    outputs(3572) <= not(layer2_outputs(3344));
    outputs(3573) <= not((layer2_outputs(6809)) xor (layer2_outputs(3615)));
    outputs(3574) <= not((layer2_outputs(8971)) xor (layer2_outputs(9717)));
    outputs(3575) <= not(layer2_outputs(7839));
    outputs(3576) <= not(layer2_outputs(7057)) or (layer2_outputs(1006));
    outputs(3577) <= not(layer2_outputs(6003));
    outputs(3578) <= layer2_outputs(8081);
    outputs(3579) <= layer2_outputs(5768);
    outputs(3580) <= layer2_outputs(6929);
    outputs(3581) <= layer2_outputs(6378);
    outputs(3582) <= (layer2_outputs(9166)) and not (layer2_outputs(2737));
    outputs(3583) <= not(layer2_outputs(769));
    outputs(3584) <= layer2_outputs(3891);
    outputs(3585) <= (layer2_outputs(3865)) and (layer2_outputs(2059));
    outputs(3586) <= not(layer2_outputs(1702)) or (layer2_outputs(7920));
    outputs(3587) <= not(layer2_outputs(5676));
    outputs(3588) <= (layer2_outputs(1147)) and (layer2_outputs(7308));
    outputs(3589) <= not(layer2_outputs(1833));
    outputs(3590) <= (layer2_outputs(5298)) xor (layer2_outputs(6225));
    outputs(3591) <= not((layer2_outputs(6257)) xor (layer2_outputs(7350)));
    outputs(3592) <= not(layer2_outputs(4762)) or (layer2_outputs(1589));
    outputs(3593) <= (layer2_outputs(2373)) and (layer2_outputs(6950));
    outputs(3594) <= not(layer2_outputs(729));
    outputs(3595) <= not(layer2_outputs(9181));
    outputs(3596) <= not(layer2_outputs(9754));
    outputs(3597) <= (layer2_outputs(4688)) xor (layer2_outputs(3364));
    outputs(3598) <= not(layer2_outputs(3570));
    outputs(3599) <= not(layer2_outputs(3422));
    outputs(3600) <= not((layer2_outputs(958)) xor (layer2_outputs(6813)));
    outputs(3601) <= not(layer2_outputs(275));
    outputs(3602) <= (layer2_outputs(8340)) and (layer2_outputs(9943));
    outputs(3603) <= not((layer2_outputs(4662)) or (layer2_outputs(6637)));
    outputs(3604) <= not(layer2_outputs(8981));
    outputs(3605) <= not((layer2_outputs(6359)) xor (layer2_outputs(2719)));
    outputs(3606) <= not(layer2_outputs(9249)) or (layer2_outputs(1370));
    outputs(3607) <= not(layer2_outputs(9198));
    outputs(3608) <= not((layer2_outputs(9077)) xor (layer2_outputs(3365)));
    outputs(3609) <= not(layer2_outputs(3114));
    outputs(3610) <= layer2_outputs(1936);
    outputs(3611) <= (layer2_outputs(1699)) xor (layer2_outputs(6807));
    outputs(3612) <= layer2_outputs(1145);
    outputs(3613) <= (layer2_outputs(8728)) and not (layer2_outputs(953));
    outputs(3614) <= not(layer2_outputs(4278));
    outputs(3615) <= (layer2_outputs(1951)) and not (layer2_outputs(5606));
    outputs(3616) <= (layer2_outputs(1858)) xor (layer2_outputs(8554));
    outputs(3617) <= layer2_outputs(6044);
    outputs(3618) <= not(layer2_outputs(6857)) or (layer2_outputs(4219));
    outputs(3619) <= layer2_outputs(9421);
    outputs(3620) <= (layer2_outputs(6697)) or (layer2_outputs(8915));
    outputs(3621) <= not(layer2_outputs(9026));
    outputs(3622) <= not(layer2_outputs(9655));
    outputs(3623) <= (layer2_outputs(1143)) or (layer2_outputs(5667));
    outputs(3624) <= not(layer2_outputs(3086));
    outputs(3625) <= (layer2_outputs(2734)) and not (layer2_outputs(9085));
    outputs(3626) <= not(layer2_outputs(3188));
    outputs(3627) <= not((layer2_outputs(7105)) xor (layer2_outputs(442)));
    outputs(3628) <= not((layer2_outputs(699)) xor (layer2_outputs(5770)));
    outputs(3629) <= not(layer2_outputs(6961));
    outputs(3630) <= not(layer2_outputs(908));
    outputs(3631) <= not((layer2_outputs(8695)) xor (layer2_outputs(4448)));
    outputs(3632) <= (layer2_outputs(9215)) xor (layer2_outputs(572));
    outputs(3633) <= layer2_outputs(927);
    outputs(3634) <= layer2_outputs(1075);
    outputs(3635) <= not((layer2_outputs(1521)) or (layer2_outputs(9007)));
    outputs(3636) <= (layer2_outputs(8265)) xor (layer2_outputs(8237));
    outputs(3637) <= layer2_outputs(4540);
    outputs(3638) <= layer2_outputs(7755);
    outputs(3639) <= layer2_outputs(5581);
    outputs(3640) <= layer2_outputs(7683);
    outputs(3641) <= (layer2_outputs(1501)) or (layer2_outputs(7709));
    outputs(3642) <= (layer2_outputs(8993)) and (layer2_outputs(2400));
    outputs(3643) <= (layer2_outputs(3877)) and (layer2_outputs(7499));
    outputs(3644) <= not(layer2_outputs(9981));
    outputs(3645) <= layer2_outputs(4096);
    outputs(3646) <= (layer2_outputs(638)) and not (layer2_outputs(8228));
    outputs(3647) <= layer2_outputs(9052);
    outputs(3648) <= layer2_outputs(6067);
    outputs(3649) <= layer2_outputs(9311);
    outputs(3650) <= not((layer2_outputs(693)) xor (layer2_outputs(6168)));
    outputs(3651) <= layer2_outputs(4821);
    outputs(3652) <= not((layer2_outputs(3914)) xor (layer2_outputs(6705)));
    outputs(3653) <= layer2_outputs(10151);
    outputs(3654) <= (layer2_outputs(8629)) and (layer2_outputs(1896));
    outputs(3655) <= not(layer2_outputs(3451));
    outputs(3656) <= not((layer2_outputs(2630)) xor (layer2_outputs(4180)));
    outputs(3657) <= not(layer2_outputs(3110));
    outputs(3658) <= (layer2_outputs(7947)) xor (layer2_outputs(3825));
    outputs(3659) <= (layer2_outputs(3580)) and not (layer2_outputs(5703));
    outputs(3660) <= not(layer2_outputs(3804));
    outputs(3661) <= not(layer2_outputs(3548));
    outputs(3662) <= not(layer2_outputs(1600));
    outputs(3663) <= (layer2_outputs(8916)) xor (layer2_outputs(9192));
    outputs(3664) <= not(layer2_outputs(552));
    outputs(3665) <= (layer2_outputs(9371)) and not (layer2_outputs(3166));
    outputs(3666) <= not(layer2_outputs(1875));
    outputs(3667) <= not((layer2_outputs(3791)) xor (layer2_outputs(3149)));
    outputs(3668) <= not(layer2_outputs(1617));
    outputs(3669) <= (layer2_outputs(144)) and not (layer2_outputs(8499));
    outputs(3670) <= not((layer2_outputs(4266)) xor (layer2_outputs(2283)));
    outputs(3671) <= layer2_outputs(1388);
    outputs(3672) <= (layer2_outputs(780)) xor (layer2_outputs(4236));
    outputs(3673) <= not(layer2_outputs(6588));
    outputs(3674) <= layer2_outputs(9014);
    outputs(3675) <= (layer2_outputs(764)) xor (layer2_outputs(3216));
    outputs(3676) <= not((layer2_outputs(6687)) and (layer2_outputs(1975)));
    outputs(3677) <= not(layer2_outputs(9304));
    outputs(3678) <= layer2_outputs(3870);
    outputs(3679) <= not(layer2_outputs(7007));
    outputs(3680) <= layer2_outputs(5451);
    outputs(3681) <= not(layer2_outputs(2933));
    outputs(3682) <= not((layer2_outputs(4615)) xor (layer2_outputs(652)));
    outputs(3683) <= layer2_outputs(9519);
    outputs(3684) <= (layer2_outputs(3783)) xor (layer2_outputs(9632));
    outputs(3685) <= not(layer2_outputs(7086));
    outputs(3686) <= not((layer2_outputs(3819)) and (layer2_outputs(1031)));
    outputs(3687) <= layer2_outputs(3175);
    outputs(3688) <= (layer2_outputs(2503)) and (layer2_outputs(5338));
    outputs(3689) <= not(layer2_outputs(9145)) or (layer2_outputs(6540));
    outputs(3690) <= not(layer2_outputs(93));
    outputs(3691) <= layer2_outputs(2905);
    outputs(3692) <= layer2_outputs(911);
    outputs(3693) <= (layer2_outputs(7368)) and (layer2_outputs(980));
    outputs(3694) <= layer2_outputs(7080);
    outputs(3695) <= not(layer2_outputs(4759));
    outputs(3696) <= (layer2_outputs(2847)) and not (layer2_outputs(4164));
    outputs(3697) <= layer2_outputs(1750);
    outputs(3698) <= layer2_outputs(1616);
    outputs(3699) <= not((layer2_outputs(9918)) xor (layer2_outputs(10070)));
    outputs(3700) <= not(layer2_outputs(8214));
    outputs(3701) <= layer2_outputs(8301);
    outputs(3702) <= (layer2_outputs(9241)) and not (layer2_outputs(3295));
    outputs(3703) <= layer2_outputs(7378);
    outputs(3704) <= layer2_outputs(7373);
    outputs(3705) <= not(layer2_outputs(1709));
    outputs(3706) <= (layer2_outputs(5977)) and not (layer2_outputs(8787));
    outputs(3707) <= not((layer2_outputs(2965)) xor (layer2_outputs(144)));
    outputs(3708) <= not((layer2_outputs(3371)) xor (layer2_outputs(2645)));
    outputs(3709) <= (layer2_outputs(7173)) xor (layer2_outputs(4206));
    outputs(3710) <= layer2_outputs(1151);
    outputs(3711) <= layer2_outputs(10118);
    outputs(3712) <= not(layer2_outputs(4826));
    outputs(3713) <= not(layer2_outputs(9330));
    outputs(3714) <= (layer2_outputs(9957)) and (layer2_outputs(2776));
    outputs(3715) <= (layer2_outputs(3262)) and (layer2_outputs(6704));
    outputs(3716) <= not(layer2_outputs(8062));
    outputs(3717) <= not(layer2_outputs(10124));
    outputs(3718) <= (layer2_outputs(6875)) xor (layer2_outputs(3212));
    outputs(3719) <= layer2_outputs(2131);
    outputs(3720) <= not((layer2_outputs(3247)) xor (layer2_outputs(5011)));
    outputs(3721) <= layer2_outputs(1177);
    outputs(3722) <= layer2_outputs(9341);
    outputs(3723) <= not(layer2_outputs(9372));
    outputs(3724) <= not(layer2_outputs(9086));
    outputs(3725) <= (layer2_outputs(3721)) or (layer2_outputs(510));
    outputs(3726) <= layer2_outputs(5325);
    outputs(3727) <= not(layer2_outputs(2021));
    outputs(3728) <= (layer2_outputs(3075)) xor (layer2_outputs(4853));
    outputs(3729) <= not(layer2_outputs(1328));
    outputs(3730) <= not(layer2_outputs(8275));
    outputs(3731) <= not((layer2_outputs(8924)) xor (layer2_outputs(10149)));
    outputs(3732) <= layer2_outputs(8912);
    outputs(3733) <= (layer2_outputs(712)) and (layer2_outputs(9499));
    outputs(3734) <= (layer2_outputs(6384)) and not (layer2_outputs(4952));
    outputs(3735) <= not(layer2_outputs(4342)) or (layer2_outputs(6750));
    outputs(3736) <= not(layer2_outputs(7932));
    outputs(3737) <= (layer2_outputs(9596)) xor (layer2_outputs(6806));
    outputs(3738) <= (layer2_outputs(1111)) and (layer2_outputs(9854));
    outputs(3739) <= not((layer2_outputs(1340)) xor (layer2_outputs(6345)));
    outputs(3740) <= layer2_outputs(2279);
    outputs(3741) <= not((layer2_outputs(585)) xor (layer2_outputs(5004)));
    outputs(3742) <= not(layer2_outputs(162));
    outputs(3743) <= not(layer2_outputs(3657));
    outputs(3744) <= not(layer2_outputs(1868));
    outputs(3745) <= (layer2_outputs(2281)) and not (layer2_outputs(6392));
    outputs(3746) <= not(layer2_outputs(2146));
    outputs(3747) <= not(layer2_outputs(7892));
    outputs(3748) <= (layer2_outputs(7787)) and (layer2_outputs(9664));
    outputs(3749) <= not(layer2_outputs(2592));
    outputs(3750) <= layer2_outputs(10042);
    outputs(3751) <= (layer2_outputs(442)) xor (layer2_outputs(1087));
    outputs(3752) <= layer2_outputs(3258);
    outputs(3753) <= not(layer2_outputs(5156));
    outputs(3754) <= not((layer2_outputs(5323)) and (layer2_outputs(506)));
    outputs(3755) <= not(layer2_outputs(2959)) or (layer2_outputs(8107));
    outputs(3756) <= not((layer2_outputs(1797)) and (layer2_outputs(9937)));
    outputs(3757) <= layer2_outputs(6974);
    outputs(3758) <= (layer2_outputs(4024)) and not (layer2_outputs(5658));
    outputs(3759) <= layer2_outputs(944);
    outputs(3760) <= not(layer2_outputs(2614));
    outputs(3761) <= not(layer2_outputs(7863)) or (layer2_outputs(6931));
    outputs(3762) <= not(layer2_outputs(736));
    outputs(3763) <= (layer2_outputs(3756)) xor (layer2_outputs(4519));
    outputs(3764) <= layer2_outputs(9766);
    outputs(3765) <= (layer2_outputs(1610)) and not (layer2_outputs(886));
    outputs(3766) <= not(layer2_outputs(6648)) or (layer2_outputs(8393));
    outputs(3767) <= not((layer2_outputs(1641)) and (layer2_outputs(5983)));
    outputs(3768) <= not(layer2_outputs(894));
    outputs(3769) <= not(layer2_outputs(5910));
    outputs(3770) <= not(layer2_outputs(5554));
    outputs(3771) <= layer2_outputs(8326);
    outputs(3772) <= not(layer2_outputs(4991));
    outputs(3773) <= (layer2_outputs(876)) and not (layer2_outputs(9403));
    outputs(3774) <= not((layer2_outputs(6436)) and (layer2_outputs(7724)));
    outputs(3775) <= (layer2_outputs(118)) or (layer2_outputs(818));
    outputs(3776) <= layer2_outputs(6000);
    outputs(3777) <= layer2_outputs(322);
    outputs(3778) <= not(layer2_outputs(740));
    outputs(3779) <= not(layer2_outputs(4225));
    outputs(3780) <= (layer2_outputs(5482)) and not (layer2_outputs(1162));
    outputs(3781) <= (layer2_outputs(218)) and not (layer2_outputs(2786));
    outputs(3782) <= (layer2_outputs(9554)) and (layer2_outputs(5534));
    outputs(3783) <= not((layer2_outputs(8087)) xor (layer2_outputs(1573)));
    outputs(3784) <= (layer2_outputs(6779)) and not (layer2_outputs(7220));
    outputs(3785) <= not(layer2_outputs(10211));
    outputs(3786) <= layer2_outputs(3770);
    outputs(3787) <= not(layer2_outputs(3946));
    outputs(3788) <= not((layer2_outputs(3988)) xor (layer2_outputs(9634)));
    outputs(3789) <= layer2_outputs(2298);
    outputs(3790) <= not((layer2_outputs(5072)) or (layer2_outputs(6888)));
    outputs(3791) <= not(layer2_outputs(5608));
    outputs(3792) <= layer2_outputs(4371);
    outputs(3793) <= (layer2_outputs(967)) and not (layer2_outputs(5067));
    outputs(3794) <= (layer2_outputs(1305)) xor (layer2_outputs(2220));
    outputs(3795) <= (layer2_outputs(3872)) and not (layer2_outputs(2939));
    outputs(3796) <= not(layer2_outputs(3495)) or (layer2_outputs(6691));
    outputs(3797) <= not(layer2_outputs(3986));
    outputs(3798) <= not(layer2_outputs(7019));
    outputs(3799) <= layer2_outputs(4804);
    outputs(3800) <= not(layer2_outputs(3439));
    outputs(3801) <= not((layer2_outputs(5060)) xor (layer2_outputs(8395)));
    outputs(3802) <= not(layer2_outputs(6641));
    outputs(3803) <= not(layer2_outputs(641));
    outputs(3804) <= layer2_outputs(8768);
    outputs(3805) <= not(layer2_outputs(9628));
    outputs(3806) <= not(layer2_outputs(1813));
    outputs(3807) <= layer2_outputs(4938);
    outputs(3808) <= not((layer2_outputs(2750)) or (layer2_outputs(686)));
    outputs(3809) <= layer2_outputs(6650);
    outputs(3810) <= not(layer2_outputs(508)) or (layer2_outputs(4506));
    outputs(3811) <= not(layer2_outputs(2455));
    outputs(3812) <= (layer2_outputs(6109)) and not (layer2_outputs(2360));
    outputs(3813) <= (layer2_outputs(6464)) and (layer2_outputs(7884));
    outputs(3814) <= not(layer2_outputs(997));
    outputs(3815) <= not(layer2_outputs(6426));
    outputs(3816) <= not(layer2_outputs(7765));
    outputs(3817) <= not(layer2_outputs(1327)) or (layer2_outputs(576));
    outputs(3818) <= (layer2_outputs(9950)) xor (layer2_outputs(269));
    outputs(3819) <= (layer2_outputs(1870)) and not (layer2_outputs(4012));
    outputs(3820) <= layer2_outputs(3018);
    outputs(3821) <= (layer2_outputs(6041)) xor (layer2_outputs(2471));
    outputs(3822) <= layer2_outputs(1382);
    outputs(3823) <= not(layer2_outputs(5732));
    outputs(3824) <= (layer2_outputs(9951)) xor (layer2_outputs(7572));
    outputs(3825) <= layer2_outputs(9546);
    outputs(3826) <= not((layer2_outputs(354)) xor (layer2_outputs(1014)));
    outputs(3827) <= not(layer2_outputs(318));
    outputs(3828) <= not((layer2_outputs(2178)) xor (layer2_outputs(4728)));
    outputs(3829) <= not(layer2_outputs(3749));
    outputs(3830) <= layer2_outputs(9409);
    outputs(3831) <= not((layer2_outputs(2758)) or (layer2_outputs(9605)));
    outputs(3832) <= layer2_outputs(1155);
    outputs(3833) <= layer2_outputs(5956);
    outputs(3834) <= (layer2_outputs(7423)) xor (layer2_outputs(1736));
    outputs(3835) <= layer2_outputs(9011);
    outputs(3836) <= not(layer2_outputs(28));
    outputs(3837) <= (layer2_outputs(8923)) and (layer2_outputs(5694));
    outputs(3838) <= (layer2_outputs(6487)) or (layer2_outputs(9815));
    outputs(3839) <= (layer2_outputs(5659)) xor (layer2_outputs(5168));
    outputs(3840) <= (layer2_outputs(7625)) and not (layer2_outputs(5834));
    outputs(3841) <= layer2_outputs(6660);
    outputs(3842) <= not(layer2_outputs(1136));
    outputs(3843) <= not(layer2_outputs(1327));
    outputs(3844) <= not(layer2_outputs(8560));
    outputs(3845) <= layer2_outputs(9237);
    outputs(3846) <= not(layer2_outputs(162));
    outputs(3847) <= layer2_outputs(5520);
    outputs(3848) <= layer2_outputs(4286);
    outputs(3849) <= not((layer2_outputs(6610)) or (layer2_outputs(2296)));
    outputs(3850) <= not(layer2_outputs(1334));
    outputs(3851) <= layer2_outputs(5384);
    outputs(3852) <= layer2_outputs(6122);
    outputs(3853) <= not(layer2_outputs(4529));
    outputs(3854) <= not((layer2_outputs(4227)) xor (layer2_outputs(1835)));
    outputs(3855) <= layer2_outputs(9449);
    outputs(3856) <= not((layer2_outputs(8941)) xor (layer2_outputs(2552)));
    outputs(3857) <= layer2_outputs(8658);
    outputs(3858) <= (layer2_outputs(323)) xor (layer2_outputs(3602));
    outputs(3859) <= not(layer2_outputs(4195));
    outputs(3860) <= not((layer2_outputs(8293)) xor (layer2_outputs(7634)));
    outputs(3861) <= not((layer2_outputs(4933)) and (layer2_outputs(255)));
    outputs(3862) <= layer2_outputs(5734);
    outputs(3863) <= layer2_outputs(6943);
    outputs(3864) <= not((layer2_outputs(9268)) or (layer2_outputs(2186)));
    outputs(3865) <= not(layer2_outputs(952));
    outputs(3866) <= not((layer2_outputs(1560)) and (layer2_outputs(8392)));
    outputs(3867) <= not(layer2_outputs(9791));
    outputs(3868) <= (layer2_outputs(7460)) xor (layer2_outputs(9973));
    outputs(3869) <= not(layer2_outputs(9522));
    outputs(3870) <= not(layer2_outputs(5157));
    outputs(3871) <= not(layer2_outputs(3608));
    outputs(3872) <= (layer2_outputs(8855)) and (layer2_outputs(6434));
    outputs(3873) <= layer2_outputs(8570);
    outputs(3874) <= not((layer2_outputs(2377)) xor (layer2_outputs(8230)));
    outputs(3875) <= not(layer2_outputs(1063));
    outputs(3876) <= (layer2_outputs(7583)) and not (layer2_outputs(590));
    outputs(3877) <= not(layer2_outputs(6106));
    outputs(3878) <= layer2_outputs(2048);
    outputs(3879) <= not(layer2_outputs(3764));
    outputs(3880) <= not(layer2_outputs(6861));
    outputs(3881) <= not(layer2_outputs(9878));
    outputs(3882) <= not(layer2_outputs(8125)) or (layer2_outputs(9776));
    outputs(3883) <= layer2_outputs(8778);
    outputs(3884) <= (layer2_outputs(3910)) and not (layer2_outputs(5152));
    outputs(3885) <= (layer2_outputs(7567)) and not (layer2_outputs(5541));
    outputs(3886) <= not(layer2_outputs(1425));
    outputs(3887) <= not((layer2_outputs(2472)) xor (layer2_outputs(4251)));
    outputs(3888) <= not(layer2_outputs(4040));
    outputs(3889) <= layer2_outputs(2577);
    outputs(3890) <= layer2_outputs(9210);
    outputs(3891) <= (layer2_outputs(1243)) xor (layer2_outputs(8140));
    outputs(3892) <= not(layer2_outputs(4171)) or (layer2_outputs(5496));
    outputs(3893) <= not(layer2_outputs(6450));
    outputs(3894) <= (layer2_outputs(6733)) and not (layer2_outputs(1765));
    outputs(3895) <= layer2_outputs(4576);
    outputs(3896) <= not(layer2_outputs(8766));
    outputs(3897) <= not(layer2_outputs(4634));
    outputs(3898) <= not(layer2_outputs(2615));
    outputs(3899) <= (layer2_outputs(1965)) xor (layer2_outputs(9146));
    outputs(3900) <= not((layer2_outputs(5565)) or (layer2_outputs(3668)));
    outputs(3901) <= not(layer2_outputs(5395));
    outputs(3902) <= (layer2_outputs(10230)) and not (layer2_outputs(3379));
    outputs(3903) <= (layer2_outputs(9336)) and not (layer2_outputs(1969));
    outputs(3904) <= layer2_outputs(9664);
    outputs(3905) <= (layer2_outputs(10106)) and (layer2_outputs(5535));
    outputs(3906) <= not(layer2_outputs(831));
    outputs(3907) <= not(layer2_outputs(2981));
    outputs(3908) <= not(layer2_outputs(5002));
    outputs(3909) <= layer2_outputs(6390);
    outputs(3910) <= (layer2_outputs(960)) xor (layer2_outputs(7695));
    outputs(3911) <= layer2_outputs(8949);
    outputs(3912) <= not(layer2_outputs(2516));
    outputs(3913) <= layer2_outputs(6360);
    outputs(3914) <= (layer2_outputs(4855)) xor (layer2_outputs(6163));
    outputs(3915) <= layer2_outputs(2099);
    outputs(3916) <= (layer2_outputs(1720)) and not (layer2_outputs(594));
    outputs(3917) <= (layer2_outputs(5698)) or (layer2_outputs(6105));
    outputs(3918) <= layer2_outputs(4620);
    outputs(3919) <= not(layer2_outputs(4326));
    outputs(3920) <= not(layer2_outputs(4748));
    outputs(3921) <= not((layer2_outputs(2425)) xor (layer2_outputs(1516)));
    outputs(3922) <= not(layer2_outputs(9741)) or (layer2_outputs(8241));
    outputs(3923) <= layer2_outputs(8189);
    outputs(3924) <= (layer2_outputs(5277)) and (layer2_outputs(9035));
    outputs(3925) <= not(layer2_outputs(8586)) or (layer2_outputs(4076));
    outputs(3926) <= (layer2_outputs(7173)) xor (layer2_outputs(6323));
    outputs(3927) <= not(layer2_outputs(1336));
    outputs(3928) <= (layer2_outputs(4838)) and not (layer2_outputs(4094));
    outputs(3929) <= (layer2_outputs(6480)) xor (layer2_outputs(7626));
    outputs(3930) <= not(layer2_outputs(3961));
    outputs(3931) <= (layer2_outputs(4152)) and not (layer2_outputs(8743));
    outputs(3932) <= (layer2_outputs(588)) or (layer2_outputs(8836));
    outputs(3933) <= (layer2_outputs(2188)) xor (layer2_outputs(8986));
    outputs(3934) <= layer2_outputs(3717);
    outputs(3935) <= not(layer2_outputs(5521));
    outputs(3936) <= (layer2_outputs(9010)) xor (layer2_outputs(4448));
    outputs(3937) <= not(layer2_outputs(1667));
    outputs(3938) <= not(layer2_outputs(8553));
    outputs(3939) <= not(layer2_outputs(3989));
    outputs(3940) <= not(layer2_outputs(7453)) or (layer2_outputs(4478));
    outputs(3941) <= not(layer2_outputs(6033)) or (layer2_outputs(1199));
    outputs(3942) <= not(layer2_outputs(8281));
    outputs(3943) <= not((layer2_outputs(8342)) or (layer2_outputs(4087)));
    outputs(3944) <= not(layer2_outputs(8204));
    outputs(3945) <= layer2_outputs(2018);
    outputs(3946) <= not((layer2_outputs(5071)) xor (layer2_outputs(2790)));
    outputs(3947) <= not(layer2_outputs(3082));
    outputs(3948) <= (layer2_outputs(6646)) or (layer2_outputs(4517));
    outputs(3949) <= (layer2_outputs(3028)) xor (layer2_outputs(4422));
    outputs(3950) <= not(layer2_outputs(5709));
    outputs(3951) <= (layer2_outputs(4811)) or (layer2_outputs(8903));
    outputs(3952) <= (layer2_outputs(4625)) xor (layer2_outputs(449));
    outputs(3953) <= not((layer2_outputs(3910)) xor (layer2_outputs(4080)));
    outputs(3954) <= (layer2_outputs(1990)) xor (layer2_outputs(7610));
    outputs(3955) <= layer2_outputs(3341);
    outputs(3956) <= not(layer2_outputs(350));
    outputs(3957) <= not((layer2_outputs(5668)) and (layer2_outputs(3358)));
    outputs(3958) <= not(layer2_outputs(1210));
    outputs(3959) <= not((layer2_outputs(2038)) xor (layer2_outputs(6375)));
    outputs(3960) <= layer2_outputs(7853);
    outputs(3961) <= layer2_outputs(957);
    outputs(3962) <= not((layer2_outputs(657)) xor (layer2_outputs(7820)));
    outputs(3963) <= not((layer2_outputs(3836)) xor (layer2_outputs(3444)));
    outputs(3964) <= not((layer2_outputs(4345)) and (layer2_outputs(1771)));
    outputs(3965) <= layer2_outputs(10125);
    outputs(3966) <= not((layer2_outputs(8536)) and (layer2_outputs(7809)));
    outputs(3967) <= not((layer2_outputs(1910)) and (layer2_outputs(3187)));
    outputs(3968) <= not((layer2_outputs(3509)) xor (layer2_outputs(2591)));
    outputs(3969) <= not(layer2_outputs(82));
    outputs(3970) <= not(layer2_outputs(172));
    outputs(3971) <= (layer2_outputs(6348)) and not (layer2_outputs(7220));
    outputs(3972) <= layer2_outputs(2166);
    outputs(3973) <= not(layer2_outputs(6295)) or (layer2_outputs(174));
    outputs(3974) <= layer2_outputs(5201);
    outputs(3975) <= not(layer2_outputs(1090));
    outputs(3976) <= (layer2_outputs(134)) and (layer2_outputs(6055));
    outputs(3977) <= (layer2_outputs(5788)) xor (layer2_outputs(4338));
    outputs(3978) <= (layer2_outputs(2057)) xor (layer2_outputs(8449));
    outputs(3979) <= not((layer2_outputs(4698)) xor (layer2_outputs(5376)));
    outputs(3980) <= not((layer2_outputs(7263)) or (layer2_outputs(4489)));
    outputs(3981) <= layer2_outputs(941);
    outputs(3982) <= (layer2_outputs(1109)) and (layer2_outputs(10203));
    outputs(3983) <= layer2_outputs(8629);
    outputs(3984) <= (layer2_outputs(7372)) and not (layer2_outputs(388));
    outputs(3985) <= layer2_outputs(6133);
    outputs(3986) <= (layer2_outputs(4375)) and not (layer2_outputs(5207));
    outputs(3987) <= layer2_outputs(3004);
    outputs(3988) <= (layer2_outputs(10129)) or (layer2_outputs(10170));
    outputs(3989) <= layer2_outputs(2234);
    outputs(3990) <= (layer2_outputs(5850)) xor (layer2_outputs(9400));
    outputs(3991) <= not((layer2_outputs(7983)) xor (layer2_outputs(4145)));
    outputs(3992) <= (layer2_outputs(375)) and not (layer2_outputs(5399));
    outputs(3993) <= not(layer2_outputs(8927));
    outputs(3994) <= not((layer2_outputs(2319)) or (layer2_outputs(3006)));
    outputs(3995) <= not(layer2_outputs(4919));
    outputs(3996) <= layer2_outputs(7260);
    outputs(3997) <= not((layer2_outputs(1171)) xor (layer2_outputs(9524)));
    outputs(3998) <= not(layer2_outputs(6778));
    outputs(3999) <= layer2_outputs(27);
    outputs(4000) <= (layer2_outputs(1734)) and (layer2_outputs(5160));
    outputs(4001) <= layer2_outputs(9725);
    outputs(4002) <= layer2_outputs(6907);
    outputs(4003) <= not((layer2_outputs(910)) or (layer2_outputs(7126)));
    outputs(4004) <= not((layer2_outputs(2495)) xor (layer2_outputs(2720)));
    outputs(4005) <= not(layer2_outputs(1981)) or (layer2_outputs(403));
    outputs(4006) <= (layer2_outputs(10006)) xor (layer2_outputs(9329));
    outputs(4007) <= not((layer2_outputs(9074)) or (layer2_outputs(328)));
    outputs(4008) <= layer2_outputs(5857);
    outputs(4009) <= layer2_outputs(8907);
    outputs(4010) <= not(layer2_outputs(3607));
    outputs(4011) <= not((layer2_outputs(2757)) xor (layer2_outputs(7119)));
    outputs(4012) <= (layer2_outputs(8875)) and not (layer2_outputs(7959));
    outputs(4013) <= not(layer2_outputs(5561));
    outputs(4014) <= layer2_outputs(10187);
    outputs(4015) <= not(layer2_outputs(8922));
    outputs(4016) <= not(layer2_outputs(511));
    outputs(4017) <= layer2_outputs(7488);
    outputs(4018) <= (layer2_outputs(8048)) and (layer2_outputs(9546));
    outputs(4019) <= layer2_outputs(2532);
    outputs(4020) <= not(layer2_outputs(9242));
    outputs(4021) <= not(layer2_outputs(2399));
    outputs(4022) <= not((layer2_outputs(119)) xor (layer2_outputs(1454)));
    outputs(4023) <= not(layer2_outputs(4694));
    outputs(4024) <= not(layer2_outputs(1085));
    outputs(4025) <= not(layer2_outputs(4837)) or (layer2_outputs(8049));
    outputs(4026) <= not(layer2_outputs(4470));
    outputs(4027) <= not((layer2_outputs(8492)) or (layer2_outputs(3800)));
    outputs(4028) <= not(layer2_outputs(2658));
    outputs(4029) <= not((layer2_outputs(9068)) xor (layer2_outputs(9370)));
    outputs(4030) <= not(layer2_outputs(5704));
    outputs(4031) <= (layer2_outputs(7543)) xor (layer2_outputs(5972));
    outputs(4032) <= (layer2_outputs(8883)) and (layer2_outputs(6607));
    outputs(4033) <= (layer2_outputs(3734)) xor (layer2_outputs(7343));
    outputs(4034) <= (layer2_outputs(6579)) xor (layer2_outputs(3662));
    outputs(4035) <= not(layer2_outputs(2093)) or (layer2_outputs(5216));
    outputs(4036) <= (layer2_outputs(7150)) xor (layer2_outputs(10035));
    outputs(4037) <= not(layer2_outputs(8800));
    outputs(4038) <= layer2_outputs(8373);
    outputs(4039) <= (layer2_outputs(6103)) xor (layer2_outputs(3507));
    outputs(4040) <= layer2_outputs(5770);
    outputs(4041) <= (layer2_outputs(1658)) xor (layer2_outputs(2366));
    outputs(4042) <= layer2_outputs(6895);
    outputs(4043) <= (layer2_outputs(4769)) xor (layer2_outputs(10201));
    outputs(4044) <= (layer2_outputs(6701)) and not (layer2_outputs(1415));
    outputs(4045) <= layer2_outputs(1427);
    outputs(4046) <= not((layer2_outputs(7529)) xor (layer2_outputs(8026)));
    outputs(4047) <= layer2_outputs(10063);
    outputs(4048) <= (layer2_outputs(6535)) and not (layer2_outputs(5136));
    outputs(4049) <= layer2_outputs(6863);
    outputs(4050) <= layer2_outputs(9045);
    outputs(4051) <= not((layer2_outputs(6784)) xor (layer2_outputs(8067)));
    outputs(4052) <= not(layer2_outputs(3103));
    outputs(4053) <= not(layer2_outputs(15)) or (layer2_outputs(3378));
    outputs(4054) <= layer2_outputs(4213);
    outputs(4055) <= (layer2_outputs(7519)) or (layer2_outputs(6113));
    outputs(4056) <= not(layer2_outputs(940));
    outputs(4057) <= not((layer2_outputs(7967)) xor (layer2_outputs(766)));
    outputs(4058) <= not(layer2_outputs(6288));
    outputs(4059) <= not(layer2_outputs(5631));
    outputs(4060) <= layer2_outputs(3529);
    outputs(4061) <= not((layer2_outputs(3549)) xor (layer2_outputs(367)));
    outputs(4062) <= (layer2_outputs(31)) xor (layer2_outputs(8206));
    outputs(4063) <= not((layer2_outputs(7542)) xor (layer2_outputs(7564)));
    outputs(4064) <= not((layer2_outputs(2886)) xor (layer2_outputs(9129)));
    outputs(4065) <= not(layer2_outputs(5793));
    outputs(4066) <= not(layer2_outputs(9572));
    outputs(4067) <= not((layer2_outputs(5167)) or (layer2_outputs(8047)));
    outputs(4068) <= (layer2_outputs(7451)) and not (layer2_outputs(2643));
    outputs(4069) <= not(layer2_outputs(7834)) or (layer2_outputs(7090));
    outputs(4070) <= not(layer2_outputs(2875));
    outputs(4071) <= (layer2_outputs(2159)) xor (layer2_outputs(4743));
    outputs(4072) <= not(layer2_outputs(9059)) or (layer2_outputs(6954));
    outputs(4073) <= layer2_outputs(2403);
    outputs(4074) <= (layer2_outputs(3850)) and (layer2_outputs(8138));
    outputs(4075) <= layer2_outputs(4371);
    outputs(4076) <= layer2_outputs(9478);
    outputs(4077) <= not((layer2_outputs(8183)) xor (layer2_outputs(3045)));
    outputs(4078) <= not(layer2_outputs(861));
    outputs(4079) <= not(layer2_outputs(3989));
    outputs(4080) <= (layer2_outputs(1468)) xor (layer2_outputs(1882));
    outputs(4081) <= not(layer2_outputs(536));
    outputs(4082) <= layer2_outputs(1958);
    outputs(4083) <= layer2_outputs(3728);
    outputs(4084) <= layer2_outputs(5622);
    outputs(4085) <= not((layer2_outputs(598)) or (layer2_outputs(3230)));
    outputs(4086) <= not((layer2_outputs(8077)) xor (layer2_outputs(9575)));
    outputs(4087) <= not(layer2_outputs(3329));
    outputs(4088) <= not(layer2_outputs(9991));
    outputs(4089) <= (layer2_outputs(4096)) and not (layer2_outputs(8816));
    outputs(4090) <= not(layer2_outputs(828));
    outputs(4091) <= (layer2_outputs(7619)) xor (layer2_outputs(5227));
    outputs(4092) <= (layer2_outputs(8561)) xor (layer2_outputs(7016));
    outputs(4093) <= not(layer2_outputs(1663));
    outputs(4094) <= not(layer2_outputs(7696));
    outputs(4095) <= not(layer2_outputs(4406));
    outputs(4096) <= not(layer2_outputs(4882));
    outputs(4097) <= not((layer2_outputs(9449)) xor (layer2_outputs(6256)));
    outputs(4098) <= not(layer2_outputs(8628)) or (layer2_outputs(9845));
    outputs(4099) <= not((layer2_outputs(1275)) xor (layer2_outputs(709)));
    outputs(4100) <= not((layer2_outputs(9718)) and (layer2_outputs(9459)));
    outputs(4101) <= not(layer2_outputs(928));
    outputs(4102) <= (layer2_outputs(1459)) and not (layer2_outputs(7346));
    outputs(4103) <= layer2_outputs(6316);
    outputs(4104) <= (layer2_outputs(6080)) or (layer2_outputs(4516));
    outputs(4105) <= not(layer2_outputs(9471));
    outputs(4106) <= not((layer2_outputs(493)) or (layer2_outputs(9106)));
    outputs(4107) <= (layer2_outputs(8246)) and not (layer2_outputs(4528));
    outputs(4108) <= not((layer2_outputs(1273)) and (layer2_outputs(5139)));
    outputs(4109) <= (layer2_outputs(8539)) and (layer2_outputs(4113));
    outputs(4110) <= layer2_outputs(1964);
    outputs(4111) <= (layer2_outputs(2880)) xor (layer2_outputs(6942));
    outputs(4112) <= layer2_outputs(7063);
    outputs(4113) <= not(layer2_outputs(3676));
    outputs(4114) <= layer2_outputs(3499);
    outputs(4115) <= layer2_outputs(6947);
    outputs(4116) <= not(layer2_outputs(6766));
    outputs(4117) <= layer2_outputs(6625);
    outputs(4118) <= layer2_outputs(4979);
    outputs(4119) <= (layer2_outputs(1508)) xor (layer2_outputs(1882));
    outputs(4120) <= not(layer2_outputs(123));
    outputs(4121) <= layer2_outputs(3009);
    outputs(4122) <= layer2_outputs(8898);
    outputs(4123) <= (layer2_outputs(937)) and (layer2_outputs(6918));
    outputs(4124) <= not(layer2_outputs(5205));
    outputs(4125) <= not(layer2_outputs(8645));
    outputs(4126) <= not(layer2_outputs(1262));
    outputs(4127) <= not(layer2_outputs(2773));
    outputs(4128) <= (layer2_outputs(6703)) and not (layer2_outputs(8643));
    outputs(4129) <= not(layer2_outputs(9368));
    outputs(4130) <= layer2_outputs(733);
    outputs(4131) <= not(layer2_outputs(2957));
    outputs(4132) <= not(layer2_outputs(7749));
    outputs(4133) <= not(layer2_outputs(1122));
    outputs(4134) <= not(layer2_outputs(7039));
    outputs(4135) <= not((layer2_outputs(176)) xor (layer2_outputs(1924)));
    outputs(4136) <= not((layer2_outputs(6257)) or (layer2_outputs(4718)));
    outputs(4137) <= layer2_outputs(1366);
    outputs(4138) <= not((layer2_outputs(7280)) xor (layer2_outputs(4856)));
    outputs(4139) <= (layer2_outputs(4982)) and not (layer2_outputs(9605));
    outputs(4140) <= layer2_outputs(3929);
    outputs(4141) <= (layer2_outputs(1670)) or (layer2_outputs(7896));
    outputs(4142) <= (layer2_outputs(9746)) and not (layer2_outputs(6282));
    outputs(4143) <= not(layer2_outputs(5584));
    outputs(4144) <= not(layer2_outputs(2833));
    outputs(4145) <= not(layer2_outputs(9801)) or (layer2_outputs(3382));
    outputs(4146) <= layer2_outputs(2222);
    outputs(4147) <= not(layer2_outputs(4934));
    outputs(4148) <= layer2_outputs(3892);
    outputs(4149) <= not(layer2_outputs(5890));
    outputs(4150) <= not((layer2_outputs(7412)) or (layer2_outputs(2677)));
    outputs(4151) <= (layer2_outputs(3083)) and (layer2_outputs(10159));
    outputs(4152) <= not((layer2_outputs(3537)) xor (layer2_outputs(2599)));
    outputs(4153) <= (layer2_outputs(7665)) or (layer2_outputs(9579));
    outputs(4154) <= layer2_outputs(10100);
    outputs(4155) <= layer2_outputs(3051);
    outputs(4156) <= (layer2_outputs(8321)) xor (layer2_outputs(5121));
    outputs(4157) <= not((layer2_outputs(2944)) or (layer2_outputs(8511)));
    outputs(4158) <= layer2_outputs(4008);
    outputs(4159) <= layer2_outputs(8635);
    outputs(4160) <= not(layer2_outputs(3980));
    outputs(4161) <= (layer2_outputs(7096)) xor (layer2_outputs(5111));
    outputs(4162) <= (layer2_outputs(6281)) xor (layer2_outputs(3323));
    outputs(4163) <= not(layer2_outputs(7992));
    outputs(4164) <= layer2_outputs(2148);
    outputs(4165) <= not(layer2_outputs(3973));
    outputs(4166) <= not(layer2_outputs(4247));
    outputs(4167) <= not(layer2_outputs(9974));
    outputs(4168) <= (layer2_outputs(8930)) and not (layer2_outputs(1402));
    outputs(4169) <= layer2_outputs(6887);
    outputs(4170) <= not(layer2_outputs(4853));
    outputs(4171) <= not((layer2_outputs(3536)) xor (layer2_outputs(9879)));
    outputs(4172) <= not(layer2_outputs(4307));
    outputs(4173) <= (layer2_outputs(9540)) and not (layer2_outputs(659));
    outputs(4174) <= not(layer2_outputs(2228));
    outputs(4175) <= not((layer2_outputs(6159)) xor (layer2_outputs(1779)));
    outputs(4176) <= (layer2_outputs(4387)) or (layer2_outputs(4318));
    outputs(4177) <= (layer2_outputs(8989)) xor (layer2_outputs(10015));
    outputs(4178) <= not((layer2_outputs(1534)) xor (layer2_outputs(1819)));
    outputs(4179) <= layer2_outputs(1233);
    outputs(4180) <= not(layer2_outputs(10183));
    outputs(4181) <= layer2_outputs(3280);
    outputs(4182) <= (layer2_outputs(235)) and not (layer2_outputs(1458));
    outputs(4183) <= not(layer2_outputs(1378));
    outputs(4184) <= layer2_outputs(2497);
    outputs(4185) <= (layer2_outputs(3654)) xor (layer2_outputs(1269));
    outputs(4186) <= (layer2_outputs(2785)) xor (layer2_outputs(6727));
    outputs(4187) <= not(layer2_outputs(5580));
    outputs(4188) <= not(layer2_outputs(9893));
    outputs(4189) <= layer2_outputs(6679);
    outputs(4190) <= layer2_outputs(7604);
    outputs(4191) <= layer2_outputs(5505);
    outputs(4192) <= not(layer2_outputs(9106));
    outputs(4193) <= not((layer2_outputs(6927)) xor (layer2_outputs(10006)));
    outputs(4194) <= not((layer2_outputs(5413)) and (layer2_outputs(6310)));
    outputs(4195) <= not(layer2_outputs(830));
    outputs(4196) <= (layer2_outputs(4582)) xor (layer2_outputs(5590));
    outputs(4197) <= layer2_outputs(6135);
    outputs(4198) <= not(layer2_outputs(7338));
    outputs(4199) <= not(layer2_outputs(5079));
    outputs(4200) <= (layer2_outputs(1682)) xor (layer2_outputs(2616));
    outputs(4201) <= not(layer2_outputs(8209));
    outputs(4202) <= not(layer2_outputs(1921));
    outputs(4203) <= not((layer2_outputs(60)) or (layer2_outputs(4642)));
    outputs(4204) <= (layer2_outputs(6049)) xor (layer2_outputs(8104));
    outputs(4205) <= layer2_outputs(4479);
    outputs(4206) <= not(layer2_outputs(1411)) or (layer2_outputs(10173));
    outputs(4207) <= not((layer2_outputs(2325)) or (layer2_outputs(3846)));
    outputs(4208) <= layer2_outputs(3014);
    outputs(4209) <= not(layer2_outputs(9639));
    outputs(4210) <= (layer2_outputs(5164)) xor (layer2_outputs(10066));
    outputs(4211) <= (layer2_outputs(2889)) xor (layer2_outputs(3037));
    outputs(4212) <= (layer2_outputs(6891)) xor (layer2_outputs(3844));
    outputs(4213) <= layer2_outputs(2946);
    outputs(4214) <= not(layer2_outputs(4255));
    outputs(4215) <= layer2_outputs(569);
    outputs(4216) <= not((layer2_outputs(1830)) xor (layer2_outputs(1)));
    outputs(4217) <= (layer2_outputs(1335)) and (layer2_outputs(4876));
    outputs(4218) <= not(layer2_outputs(8445));
    outputs(4219) <= not((layer2_outputs(5523)) xor (layer2_outputs(7288)));
    outputs(4220) <= not((layer2_outputs(6517)) and (layer2_outputs(7755)));
    outputs(4221) <= not((layer2_outputs(9361)) xor (layer2_outputs(10126)));
    outputs(4222) <= layer2_outputs(5053);
    outputs(4223) <= not(layer2_outputs(10184));
    outputs(4224) <= layer2_outputs(8380);
    outputs(4225) <= not(layer2_outputs(4212));
    outputs(4226) <= layer2_outputs(970);
    outputs(4227) <= layer2_outputs(4238);
    outputs(4228) <= not(layer2_outputs(5331)) or (layer2_outputs(3280));
    outputs(4229) <= not((layer2_outputs(8820)) xor (layer2_outputs(250)));
    outputs(4230) <= not(layer2_outputs(3419));
    outputs(4231) <= not(layer2_outputs(5203)) or (layer2_outputs(5621));
    outputs(4232) <= not(layer2_outputs(9549));
    outputs(4233) <= (layer2_outputs(4867)) and not (layer2_outputs(10031));
    outputs(4234) <= layer2_outputs(8123);
    outputs(4235) <= not(layer2_outputs(875)) or (layer2_outputs(10134));
    outputs(4236) <= not(layer2_outputs(7786));
    outputs(4237) <= layer2_outputs(6251);
    outputs(4238) <= not(layer2_outputs(8976));
    outputs(4239) <= layer2_outputs(9291);
    outputs(4240) <= not(layer2_outputs(9324));
    outputs(4241) <= layer2_outputs(9349);
    outputs(4242) <= not(layer2_outputs(1998));
    outputs(4243) <= layer2_outputs(8017);
    outputs(4244) <= not((layer2_outputs(1131)) or (layer2_outputs(666)));
    outputs(4245) <= (layer2_outputs(7816)) and not (layer2_outputs(5718));
    outputs(4246) <= not(layer2_outputs(1171)) or (layer2_outputs(4357));
    outputs(4247) <= not(layer2_outputs(5482));
    outputs(4248) <= not(layer2_outputs(4846));
    outputs(4249) <= layer2_outputs(1928);
    outputs(4250) <= (layer2_outputs(9034)) or (layer2_outputs(10137));
    outputs(4251) <= not(layer2_outputs(7378));
    outputs(4252) <= (layer2_outputs(6887)) and not (layer2_outputs(9686));
    outputs(4253) <= layer2_outputs(9507);
    outputs(4254) <= not((layer2_outputs(82)) xor (layer2_outputs(4171)));
    outputs(4255) <= layer2_outputs(4074);
    outputs(4256) <= (layer2_outputs(2739)) xor (layer2_outputs(3440));
    outputs(4257) <= not(layer2_outputs(7958)) or (layer2_outputs(4203));
    outputs(4258) <= not(layer2_outputs(4794));
    outputs(4259) <= not(layer2_outputs(4944));
    outputs(4260) <= not(layer2_outputs(1050));
    outputs(4261) <= not(layer2_outputs(3725));
    outputs(4262) <= not(layer2_outputs(3930));
    outputs(4263) <= not(layer2_outputs(292));
    outputs(4264) <= layer2_outputs(678);
    outputs(4265) <= not(layer2_outputs(8581));
    outputs(4266) <= (layer2_outputs(4815)) xor (layer2_outputs(6130));
    outputs(4267) <= not(layer2_outputs(2674));
    outputs(4268) <= layer2_outputs(2258);
    outputs(4269) <= not((layer2_outputs(1971)) and (layer2_outputs(5037)));
    outputs(4270) <= not((layer2_outputs(9021)) or (layer2_outputs(8019)));
    outputs(4271) <= not(layer2_outputs(4337));
    outputs(4272) <= layer2_outputs(7659);
    outputs(4273) <= not(layer2_outputs(6574));
    outputs(4274) <= not(layer2_outputs(5838)) or (layer2_outputs(3596));
    outputs(4275) <= not(layer2_outputs(5963));
    outputs(4276) <= layer2_outputs(8118);
    outputs(4277) <= not((layer2_outputs(4359)) xor (layer2_outputs(2484)));
    outputs(4278) <= (layer2_outputs(3105)) and not (layer2_outputs(4705));
    outputs(4279) <= not((layer2_outputs(8758)) xor (layer2_outputs(8777)));
    outputs(4280) <= layer2_outputs(1546);
    outputs(4281) <= not(layer2_outputs(4354));
    outputs(4282) <= not(layer2_outputs(2677));
    outputs(4283) <= (layer2_outputs(3987)) and not (layer2_outputs(9837));
    outputs(4284) <= not((layer2_outputs(9267)) xor (layer2_outputs(5186)));
    outputs(4285) <= layer2_outputs(8814);
    outputs(4286) <= not(layer2_outputs(8436));
    outputs(4287) <= (layer2_outputs(4218)) xor (layer2_outputs(2481));
    outputs(4288) <= (layer2_outputs(6269)) and not (layer2_outputs(6654));
    outputs(4289) <= layer2_outputs(4284);
    outputs(4290) <= (layer2_outputs(7807)) and not (layer2_outputs(1538));
    outputs(4291) <= layer2_outputs(555);
    outputs(4292) <= layer2_outputs(6604);
    outputs(4293) <= not(layer2_outputs(7468)) or (layer2_outputs(4614));
    outputs(4294) <= layer2_outputs(28);
    outputs(4295) <= not(layer2_outputs(5655));
    outputs(4296) <= not(layer2_outputs(8847));
    outputs(4297) <= not(layer2_outputs(359)) or (layer2_outputs(8894));
    outputs(4298) <= not(layer2_outputs(813));
    outputs(4299) <= not(layer2_outputs(10058));
    outputs(4300) <= (layer2_outputs(8280)) xor (layer2_outputs(5292));
    outputs(4301) <= not(layer2_outputs(1039));
    outputs(4302) <= not(layer2_outputs(9523));
    outputs(4303) <= (layer2_outputs(288)) and not (layer2_outputs(5823));
    outputs(4304) <= not(layer2_outputs(9812));
    outputs(4305) <= not(layer2_outputs(4063));
    outputs(4306) <= (layer2_outputs(4443)) or (layer2_outputs(5719));
    outputs(4307) <= (layer2_outputs(2052)) and not (layer2_outputs(6510));
    outputs(4308) <= layer2_outputs(3881);
    outputs(4309) <= not(layer2_outputs(4440)) or (layer2_outputs(3152));
    outputs(4310) <= not((layer2_outputs(5007)) and (layer2_outputs(4038)));
    outputs(4311) <= layer2_outputs(2130);
    outputs(4312) <= not((layer2_outputs(6118)) xor (layer2_outputs(3493)));
    outputs(4313) <= (layer2_outputs(3174)) xor (layer2_outputs(2407));
    outputs(4314) <= not(layer2_outputs(1786));
    outputs(4315) <= (layer2_outputs(345)) xor (layer2_outputs(56));
    outputs(4316) <= not(layer2_outputs(8929));
    outputs(4317) <= not(layer2_outputs(4438)) or (layer2_outputs(7188));
    outputs(4318) <= layer2_outputs(418);
    outputs(4319) <= not((layer2_outputs(896)) and (layer2_outputs(4329)));
    outputs(4320) <= not(layer2_outputs(7021));
    outputs(4321) <= not(layer2_outputs(8578));
    outputs(4322) <= (layer2_outputs(10002)) xor (layer2_outputs(526));
    outputs(4323) <= layer2_outputs(1946);
    outputs(4324) <= not(layer2_outputs(3884)) or (layer2_outputs(7620));
    outputs(4325) <= (layer2_outputs(3532)) xor (layer2_outputs(7123));
    outputs(4326) <= layer2_outputs(3115);
    outputs(4327) <= not(layer2_outputs(1852)) or (layer2_outputs(10011));
    outputs(4328) <= not(layer2_outputs(6332));
    outputs(4329) <= layer2_outputs(1423);
    outputs(4330) <= (layer2_outputs(4340)) xor (layer2_outputs(10140));
    outputs(4331) <= (layer2_outputs(396)) and not (layer2_outputs(5354));
    outputs(4332) <= (layer2_outputs(1191)) and (layer2_outputs(7803));
    outputs(4333) <= layer2_outputs(509);
    outputs(4334) <= layer2_outputs(181);
    outputs(4335) <= (layer2_outputs(7698)) xor (layer2_outputs(1260));
    outputs(4336) <= not(layer2_outputs(3054));
    outputs(4337) <= layer2_outputs(7218);
    outputs(4338) <= (layer2_outputs(3127)) and not (layer2_outputs(8292));
    outputs(4339) <= not(layer2_outputs(3937));
    outputs(4340) <= not((layer2_outputs(1367)) xor (layer2_outputs(3573)));
    outputs(4341) <= not((layer2_outputs(3283)) or (layer2_outputs(1043)));
    outputs(4342) <= not(layer2_outputs(6226));
    outputs(4343) <= not(layer2_outputs(7217));
    outputs(4344) <= not((layer2_outputs(7711)) and (layer2_outputs(110)));
    outputs(4345) <= (layer2_outputs(5760)) xor (layer2_outputs(5582));
    outputs(4346) <= layer2_outputs(3122);
    outputs(4347) <= (layer2_outputs(3333)) xor (layer2_outputs(7673));
    outputs(4348) <= (layer2_outputs(4414)) and not (layer2_outputs(5303));
    outputs(4349) <= not((layer2_outputs(6420)) or (layer2_outputs(2669)));
    outputs(4350) <= not((layer2_outputs(1330)) xor (layer2_outputs(717)));
    outputs(4351) <= not((layer2_outputs(5927)) or (layer2_outputs(1126)));
    outputs(4352) <= layer2_outputs(3323);
    outputs(4353) <= layer2_outputs(2250);
    outputs(4354) <= not(layer2_outputs(8201));
    outputs(4355) <= not(layer2_outputs(2568));
    outputs(4356) <= not((layer2_outputs(1203)) and (layer2_outputs(8977)));
    outputs(4357) <= layer2_outputs(9038);
    outputs(4358) <= layer2_outputs(245);
    outputs(4359) <= not(layer2_outputs(9346));
    outputs(4360) <= not(layer2_outputs(6371));
    outputs(4361) <= not((layer2_outputs(6873)) xor (layer2_outputs(7662)));
    outputs(4362) <= not(layer2_outputs(7021));
    outputs(4363) <= layer2_outputs(1176);
    outputs(4364) <= not((layer2_outputs(5726)) xor (layer2_outputs(10046)));
    outputs(4365) <= layer2_outputs(8156);
    outputs(4366) <= layer2_outputs(1077);
    outputs(4367) <= not(layer2_outputs(9617));
    outputs(4368) <= not(layer2_outputs(3737));
    outputs(4369) <= layer2_outputs(4978);
    outputs(4370) <= not((layer2_outputs(2810)) xor (layer2_outputs(7629)));
    outputs(4371) <= (layer2_outputs(8818)) or (layer2_outputs(9428));
    outputs(4372) <= layer2_outputs(3813);
    outputs(4373) <= layer2_outputs(9622);
    outputs(4374) <= not(layer2_outputs(644));
    outputs(4375) <= not(layer2_outputs(705));
    outputs(4376) <= not(layer2_outputs(7584)) or (layer2_outputs(4685));
    outputs(4377) <= not(layer2_outputs(5883));
    outputs(4378) <= (layer2_outputs(9995)) and not (layer2_outputs(2923));
    outputs(4379) <= not(layer2_outputs(6692));
    outputs(4380) <= layer2_outputs(7105);
    outputs(4381) <= not(layer2_outputs(2732));
    outputs(4382) <= (layer2_outputs(1801)) and (layer2_outputs(6186));
    outputs(4383) <= layer2_outputs(2463);
    outputs(4384) <= layer2_outputs(8402);
    outputs(4385) <= (layer2_outputs(998)) xor (layer2_outputs(8186));
    outputs(4386) <= not(layer2_outputs(8654));
    outputs(4387) <= not(layer2_outputs(5165));
    outputs(4388) <= not(layer2_outputs(1575));
    outputs(4389) <= layer2_outputs(7410);
    outputs(4390) <= not(layer2_outputs(7437));
    outputs(4391) <= not(layer2_outputs(184));
    outputs(4392) <= layer2_outputs(1490);
    outputs(4393) <= (layer2_outputs(8119)) and not (layer2_outputs(6658));
    outputs(4394) <= layer2_outputs(7410);
    outputs(4395) <= not(layer2_outputs(3776));
    outputs(4396) <= not((layer2_outputs(2321)) or (layer2_outputs(1921)));
    outputs(4397) <= (layer2_outputs(2919)) and not (layer2_outputs(4681));
    outputs(4398) <= layer2_outputs(7942);
    outputs(4399) <= not(layer2_outputs(5348)) or (layer2_outputs(7367));
    outputs(4400) <= '0';
    outputs(4401) <= layer2_outputs(6800);
    outputs(4402) <= (layer2_outputs(6203)) xor (layer2_outputs(6758));
    outputs(4403) <= (layer2_outputs(981)) and not (layer2_outputs(157));
    outputs(4404) <= layer2_outputs(5788);
    outputs(4405) <= layer2_outputs(3128);
    outputs(4406) <= layer2_outputs(3860);
    outputs(4407) <= (layer2_outputs(7973)) and (layer2_outputs(4951));
    outputs(4408) <= (layer2_outputs(2006)) xor (layer2_outputs(2884));
    outputs(4409) <= layer2_outputs(1226);
    outputs(4410) <= layer2_outputs(8824);
    outputs(4411) <= layer2_outputs(4443);
    outputs(4412) <= (layer2_outputs(5649)) and (layer2_outputs(9866));
    outputs(4413) <= not(layer2_outputs(4058)) or (layer2_outputs(618));
    outputs(4414) <= layer2_outputs(7011);
    outputs(4415) <= layer2_outputs(7598);
    outputs(4416) <= not(layer2_outputs(4666));
    outputs(4417) <= (layer2_outputs(1357)) and not (layer2_outputs(7340));
    outputs(4418) <= not(layer2_outputs(5470));
    outputs(4419) <= layer2_outputs(3251);
    outputs(4420) <= (layer2_outputs(7959)) or (layer2_outputs(684));
    outputs(4421) <= not((layer2_outputs(3568)) or (layer2_outputs(5305)));
    outputs(4422) <= layer2_outputs(5001);
    outputs(4423) <= not(layer2_outputs(8137)) or (layer2_outputs(4407));
    outputs(4424) <= (layer2_outputs(3739)) or (layer2_outputs(648));
    outputs(4425) <= layer2_outputs(6878);
    outputs(4426) <= (layer2_outputs(2670)) xor (layer2_outputs(887));
    outputs(4427) <= (layer2_outputs(2129)) and not (layer2_outputs(7599));
    outputs(4428) <= not((layer2_outputs(3650)) or (layer2_outputs(605)));
    outputs(4429) <= layer2_outputs(684);
    outputs(4430) <= not(layer2_outputs(9195));
    outputs(4431) <= layer2_outputs(8966);
    outputs(4432) <= layer2_outputs(4638);
    outputs(4433) <= (layer2_outputs(3525)) or (layer2_outputs(9497));
    outputs(4434) <= not(layer2_outputs(2320));
    outputs(4435) <= (layer2_outputs(2265)) and not (layer2_outputs(4256));
    outputs(4436) <= not(layer2_outputs(2533));
    outputs(4437) <= not((layer2_outputs(8660)) xor (layer2_outputs(6614)));
    outputs(4438) <= (layer2_outputs(5703)) xor (layer2_outputs(6108));
    outputs(4439) <= layer2_outputs(2109);
    outputs(4440) <= not((layer2_outputs(884)) xor (layer2_outputs(7465)));
    outputs(4441) <= not(layer2_outputs(3765));
    outputs(4442) <= not(layer2_outputs(8404));
    outputs(4443) <= not(layer2_outputs(7911));
    outputs(4444) <= not(layer2_outputs(231));
    outputs(4445) <= (layer2_outputs(3451)) and not (layer2_outputs(4305));
    outputs(4446) <= not(layer2_outputs(6736));
    outputs(4447) <= not((layer2_outputs(7443)) xor (layer2_outputs(7116)));
    outputs(4448) <= (layer2_outputs(7450)) and not (layer2_outputs(4686));
    outputs(4449) <= not(layer2_outputs(99));
    outputs(4450) <= not(layer2_outputs(3534)) or (layer2_outputs(1832));
    outputs(4451) <= not((layer2_outputs(9072)) and (layer2_outputs(7458)));
    outputs(4452) <= not((layer2_outputs(1631)) xor (layer2_outputs(6012)));
    outputs(4453) <= not((layer2_outputs(6222)) xor (layer2_outputs(5353)));
    outputs(4454) <= not(layer2_outputs(9288));
    outputs(4455) <= not(layer2_outputs(8098));
    outputs(4456) <= layer2_outputs(4520);
    outputs(4457) <= (layer2_outputs(5106)) xor (layer2_outputs(6069));
    outputs(4458) <= layer2_outputs(7459);
    outputs(4459) <= layer2_outputs(6117);
    outputs(4460) <= layer2_outputs(9647);
    outputs(4461) <= layer2_outputs(3467);
    outputs(4462) <= not(layer2_outputs(10192));
    outputs(4463) <= (layer2_outputs(2017)) and not (layer2_outputs(5091));
    outputs(4464) <= not(layer2_outputs(2087));
    outputs(4465) <= layer2_outputs(223);
    outputs(4466) <= layer2_outputs(9323);
    outputs(4467) <= layer2_outputs(4932);
    outputs(4468) <= (layer2_outputs(7097)) and not (layer2_outputs(9598));
    outputs(4469) <= not(layer2_outputs(8653));
    outputs(4470) <= not(layer2_outputs(9932));
    outputs(4471) <= (layer2_outputs(6971)) and not (layer2_outputs(9476));
    outputs(4472) <= (layer2_outputs(9708)) xor (layer2_outputs(9782));
    outputs(4473) <= not(layer2_outputs(3711));
    outputs(4474) <= not((layer2_outputs(3784)) or (layer2_outputs(2940)));
    outputs(4475) <= (layer2_outputs(10078)) xor (layer2_outputs(4538));
    outputs(4476) <= (layer2_outputs(9396)) and (layer2_outputs(9758));
    outputs(4477) <= layer2_outputs(7036);
    outputs(4478) <= (layer2_outputs(5911)) and not (layer2_outputs(5201));
    outputs(4479) <= not((layer2_outputs(1932)) xor (layer2_outputs(2071)));
    outputs(4480) <= not(layer2_outputs(2433));
    outputs(4481) <= (layer2_outputs(10214)) xor (layer2_outputs(9739));
    outputs(4482) <= layer2_outputs(4237);
    outputs(4483) <= layer2_outputs(409);
    outputs(4484) <= not(layer2_outputs(2162));
    outputs(4485) <= layer2_outputs(9039);
    outputs(4486) <= layer2_outputs(2223);
    outputs(4487) <= layer2_outputs(4999);
    outputs(4488) <= not((layer2_outputs(9637)) or (layer2_outputs(317)));
    outputs(4489) <= not(layer2_outputs(4549));
    outputs(4490) <= not(layer2_outputs(421));
    outputs(4491) <= not(layer2_outputs(4099));
    outputs(4492) <= not((layer2_outputs(8347)) xor (layer2_outputs(10109)));
    outputs(4493) <= not(layer2_outputs(7940));
    outputs(4494) <= layer2_outputs(7831);
    outputs(4495) <= (layer2_outputs(6388)) and not (layer2_outputs(7523));
    outputs(4496) <= (layer2_outputs(9656)) and (layer2_outputs(548));
    outputs(4497) <= (layer2_outputs(3361)) xor (layer2_outputs(2600));
    outputs(4498) <= layer2_outputs(6286);
    outputs(4499) <= (layer2_outputs(9192)) or (layer2_outputs(5628));
    outputs(4500) <= not(layer2_outputs(1271));
    outputs(4501) <= not((layer2_outputs(9047)) and (layer2_outputs(5279)));
    outputs(4502) <= not(layer2_outputs(5052));
    outputs(4503) <= (layer2_outputs(9244)) xor (layer2_outputs(4272));
    outputs(4504) <= layer2_outputs(8577);
    outputs(4505) <= (layer2_outputs(7472)) and not (layer2_outputs(6416));
    outputs(4506) <= layer2_outputs(6880);
    outputs(4507) <= not((layer2_outputs(3934)) or (layer2_outputs(5600)));
    outputs(4508) <= (layer2_outputs(7135)) and not (layer2_outputs(4254));
    outputs(4509) <= (layer2_outputs(10178)) xor (layer2_outputs(3843));
    outputs(4510) <= not(layer2_outputs(7046));
    outputs(4511) <= not(layer2_outputs(3420));
    outputs(4512) <= not((layer2_outputs(8912)) and (layer2_outputs(4628)));
    outputs(4513) <= layer2_outputs(6432);
    outputs(4514) <= (layer2_outputs(5663)) xor (layer2_outputs(7205));
    outputs(4515) <= layer2_outputs(1883);
    outputs(4516) <= not(layer2_outputs(5056)) or (layer2_outputs(1982));
    outputs(4517) <= layer2_outputs(8294);
    outputs(4518) <= (layer2_outputs(3220)) or (layer2_outputs(5352));
    outputs(4519) <= layer2_outputs(404);
    outputs(4520) <= not(layer2_outputs(2487));
    outputs(4521) <= not(layer2_outputs(3332));
    outputs(4522) <= not(layer2_outputs(4861));
    outputs(4523) <= layer2_outputs(4651);
    outputs(4524) <= layer2_outputs(3191);
    outputs(4525) <= not((layer2_outputs(9591)) xor (layer2_outputs(657)));
    outputs(4526) <= layer2_outputs(3095);
    outputs(4527) <= not((layer2_outputs(4034)) or (layer2_outputs(5418)));
    outputs(4528) <= layer2_outputs(2912);
    outputs(4529) <= (layer2_outputs(8986)) xor (layer2_outputs(8950));
    outputs(4530) <= not(layer2_outputs(9563));
    outputs(4531) <= not((layer2_outputs(6007)) xor (layer2_outputs(6523)));
    outputs(4532) <= not(layer2_outputs(2373));
    outputs(4533) <= not(layer2_outputs(8190)) or (layer2_outputs(1289));
    outputs(4534) <= (layer2_outputs(6931)) xor (layer2_outputs(386));
    outputs(4535) <= not(layer2_outputs(7114));
    outputs(4536) <= not(layer2_outputs(8946));
    outputs(4537) <= (layer2_outputs(3513)) xor (layer2_outputs(3027));
    outputs(4538) <= not(layer2_outputs(6497));
    outputs(4539) <= (layer2_outputs(8580)) and (layer2_outputs(2646));
    outputs(4540) <= not((layer2_outputs(595)) xor (layer2_outputs(4265)));
    outputs(4541) <= (layer2_outputs(192)) xor (layer2_outputs(9588));
    outputs(4542) <= not(layer2_outputs(565));
    outputs(4543) <= (layer2_outputs(6546)) and not (layer2_outputs(3417));
    outputs(4544) <= not(layer2_outputs(9941));
    outputs(4545) <= layer2_outputs(668);
    outputs(4546) <= (layer2_outputs(8076)) and (layer2_outputs(867));
    outputs(4547) <= (layer2_outputs(4493)) and not (layer2_outputs(5524));
    outputs(4548) <= not(layer2_outputs(3205));
    outputs(4549) <= layer2_outputs(2105);
    outputs(4550) <= not((layer2_outputs(2675)) or (layer2_outputs(5282)));
    outputs(4551) <= layer2_outputs(4845);
    outputs(4552) <= (layer2_outputs(9506)) xor (layer2_outputs(3349));
    outputs(4553) <= not((layer2_outputs(198)) or (layer2_outputs(8656)));
    outputs(4554) <= not((layer2_outputs(8552)) xor (layer2_outputs(3707)));
    outputs(4555) <= layer2_outputs(34);
    outputs(4556) <= (layer2_outputs(7181)) and not (layer2_outputs(9836));
    outputs(4557) <= layer2_outputs(1689);
    outputs(4558) <= layer2_outputs(9348);
    outputs(4559) <= layer2_outputs(4495);
    outputs(4560) <= not(layer2_outputs(4937));
    outputs(4561) <= (layer2_outputs(254)) and (layer2_outputs(8041));
    outputs(4562) <= not(layer2_outputs(1723));
    outputs(4563) <= (layer2_outputs(3902)) and (layer2_outputs(4747));
    outputs(4564) <= (layer2_outputs(2594)) xor (layer2_outputs(6755));
    outputs(4565) <= not(layer2_outputs(2458));
    outputs(4566) <= (layer2_outputs(2239)) and not (layer2_outputs(6102));
    outputs(4567) <= not(layer2_outputs(8352));
    outputs(4568) <= layer2_outputs(2488);
    outputs(4569) <= not(layer2_outputs(332));
    outputs(4570) <= not(layer2_outputs(7385));
    outputs(4571) <= (layer2_outputs(7978)) and not (layer2_outputs(8223));
    outputs(4572) <= layer2_outputs(8147);
    outputs(4573) <= not(layer2_outputs(227));
    outputs(4574) <= layer2_outputs(5774);
    outputs(4575) <= not((layer2_outputs(813)) or (layer2_outputs(7437)));
    outputs(4576) <= layer2_outputs(9648);
    outputs(4577) <= not(layer2_outputs(1110));
    outputs(4578) <= (layer2_outputs(692)) xor (layer2_outputs(1164));
    outputs(4579) <= layer2_outputs(8896);
    outputs(4580) <= not(layer2_outputs(5085));
    outputs(4581) <= layer2_outputs(3091);
    outputs(4582) <= layer2_outputs(6463);
    outputs(4583) <= not(layer2_outputs(8092));
    outputs(4584) <= not(layer2_outputs(8239)) or (layer2_outputs(6065));
    outputs(4585) <= (layer2_outputs(1046)) xor (layer2_outputs(1854));
    outputs(4586) <= not((layer2_outputs(8491)) or (layer2_outputs(2675)));
    outputs(4587) <= layer2_outputs(9810);
    outputs(4588) <= not((layer2_outputs(3148)) and (layer2_outputs(6511)));
    outputs(4589) <= layer2_outputs(3950);
    outputs(4590) <= (layer2_outputs(5557)) and not (layer2_outputs(10102));
    outputs(4591) <= layer2_outputs(6201);
    outputs(4592) <= not(layer2_outputs(2550));
    outputs(4593) <= not(layer2_outputs(1687)) or (layer2_outputs(10051));
    outputs(4594) <= not((layer2_outputs(6364)) xor (layer2_outputs(4668)));
    outputs(4595) <= not(layer2_outputs(9442));
    outputs(4596) <= not(layer2_outputs(3675));
    outputs(4597) <= (layer2_outputs(5713)) and not (layer2_outputs(9217));
    outputs(4598) <= (layer2_outputs(9969)) xor (layer2_outputs(9490));
    outputs(4599) <= not(layer2_outputs(4838));
    outputs(4600) <= (layer2_outputs(4318)) or (layer2_outputs(1631));
    outputs(4601) <= not(layer2_outputs(1055));
    outputs(4602) <= layer2_outputs(7864);
    outputs(4603) <= layer2_outputs(1476);
    outputs(4604) <= not((layer2_outputs(849)) xor (layer2_outputs(5961)));
    outputs(4605) <= not(layer2_outputs(1492));
    outputs(4606) <= not(layer2_outputs(2229));
    outputs(4607) <= layer2_outputs(6899);
    outputs(4608) <= not((layer2_outputs(5119)) xor (layer2_outputs(9389)));
    outputs(4609) <= not((layer2_outputs(3526)) or (layer2_outputs(1463)));
    outputs(4610) <= not(layer2_outputs(1400));
    outputs(4611) <= (layer2_outputs(9753)) and not (layer2_outputs(8352));
    outputs(4612) <= not(layer2_outputs(3476));
    outputs(4613) <= not((layer2_outputs(2832)) xor (layer2_outputs(1471)));
    outputs(4614) <= not(layer2_outputs(2787));
    outputs(4615) <= not(layer2_outputs(381));
    outputs(4616) <= not(layer2_outputs(6305));
    outputs(4617) <= not(layer2_outputs(8346));
    outputs(4618) <= not((layer2_outputs(1377)) and (layer2_outputs(5980)));
    outputs(4619) <= layer2_outputs(1077);
    outputs(4620) <= (layer2_outputs(5145)) xor (layer2_outputs(5826));
    outputs(4621) <= layer2_outputs(4664);
    outputs(4622) <= not(layer2_outputs(1076));
    outputs(4623) <= not((layer2_outputs(6587)) or (layer2_outputs(7402)));
    outputs(4624) <= layer2_outputs(2323);
    outputs(4625) <= layer2_outputs(2796);
    outputs(4626) <= layer2_outputs(458);
    outputs(4627) <= layer2_outputs(42);
    outputs(4628) <= not((layer2_outputs(5854)) xor (layer2_outputs(3810)));
    outputs(4629) <= not((layer2_outputs(6034)) or (layer2_outputs(7768)));
    outputs(4630) <= not((layer2_outputs(8631)) and (layer2_outputs(7284)));
    outputs(4631) <= (layer2_outputs(5465)) and (layer2_outputs(2446));
    outputs(4632) <= layer2_outputs(4576);
    outputs(4633) <= (layer2_outputs(2398)) xor (layer2_outputs(2672));
    outputs(4634) <= layer2_outputs(9779);
    outputs(4635) <= not((layer2_outputs(4785)) or (layer2_outputs(1045)));
    outputs(4636) <= (layer2_outputs(4424)) xor (layer2_outputs(6382));
    outputs(4637) <= layer2_outputs(6072);
    outputs(4638) <= not(layer2_outputs(10053));
    outputs(4639) <= layer2_outputs(318);
    outputs(4640) <= not(layer2_outputs(1402)) or (layer2_outputs(1614));
    outputs(4641) <= not((layer2_outputs(6943)) or (layer2_outputs(9846)));
    outputs(4642) <= not((layer2_outputs(7356)) xor (layer2_outputs(3080)));
    outputs(4643) <= not(layer2_outputs(6557));
    outputs(4644) <= not(layer2_outputs(5500));
    outputs(4645) <= (layer2_outputs(46)) xor (layer2_outputs(7701));
    outputs(4646) <= (layer2_outputs(7571)) xor (layer2_outputs(7379));
    outputs(4647) <= not(layer2_outputs(2515));
    outputs(4648) <= layer2_outputs(9213);
    outputs(4649) <= not(layer2_outputs(8396));
    outputs(4650) <= layer2_outputs(1514);
    outputs(4651) <= not(layer2_outputs(3224));
    outputs(4652) <= not(layer2_outputs(1316)) or (layer2_outputs(5069));
    outputs(4653) <= layer2_outputs(2371);
    outputs(4654) <= (layer2_outputs(5539)) and not (layer2_outputs(4603));
    outputs(4655) <= (layer2_outputs(7536)) xor (layer2_outputs(7115));
    outputs(4656) <= layer2_outputs(515);
    outputs(4657) <= layer2_outputs(8541);
    outputs(4658) <= layer2_outputs(3317);
    outputs(4659) <= not(layer2_outputs(4169));
    outputs(4660) <= (layer2_outputs(8580)) xor (layer2_outputs(1249));
    outputs(4661) <= not(layer2_outputs(9307));
    outputs(4662) <= (layer2_outputs(4319)) or (layer2_outputs(133));
    outputs(4663) <= not((layer2_outputs(4575)) xor (layer2_outputs(6009)));
    outputs(4664) <= (layer2_outputs(8879)) xor (layer2_outputs(4093));
    outputs(4665) <= layer2_outputs(9990);
    outputs(4666) <= not((layer2_outputs(4555)) or (layer2_outputs(484)));
    outputs(4667) <= layer2_outputs(7183);
    outputs(4668) <= layer2_outputs(6322);
    outputs(4669) <= (layer2_outputs(1799)) and (layer2_outputs(402));
    outputs(4670) <= layer2_outputs(3667);
    outputs(4671) <= not(layer2_outputs(9264));
    outputs(4672) <= layer2_outputs(4050);
    outputs(4673) <= layer2_outputs(5064);
    outputs(4674) <= not(layer2_outputs(6552));
    outputs(4675) <= (layer2_outputs(374)) or (layer2_outputs(8119));
    outputs(4676) <= not(layer2_outputs(3348));
    outputs(4677) <= not(layer2_outputs(5732));
    outputs(4678) <= (layer2_outputs(9788)) xor (layer2_outputs(6276));
    outputs(4679) <= not(layer2_outputs(5025));
    outputs(4680) <= (layer2_outputs(4992)) and not (layer2_outputs(5747));
    outputs(4681) <= not(layer2_outputs(369));
    outputs(4682) <= not((layer2_outputs(3346)) xor (layer2_outputs(121)));
    outputs(4683) <= not((layer2_outputs(1457)) xor (layer2_outputs(7277)));
    outputs(4684) <= not((layer2_outputs(9919)) xor (layer2_outputs(7629)));
    outputs(4685) <= layer2_outputs(9381);
    outputs(4686) <= not((layer2_outputs(5510)) xor (layer2_outputs(1906)));
    outputs(4687) <= layer2_outputs(7748);
    outputs(4688) <= not(layer2_outputs(3199));
    outputs(4689) <= layer2_outputs(10116);
    outputs(4690) <= not((layer2_outputs(1156)) xor (layer2_outputs(7227)));
    outputs(4691) <= layer2_outputs(9351);
    outputs(4692) <= not(layer2_outputs(5066)) or (layer2_outputs(7407));
    outputs(4693) <= not(layer2_outputs(4926));
    outputs(4694) <= not(layer2_outputs(4260));
    outputs(4695) <= not((layer2_outputs(2830)) and (layer2_outputs(9195)));
    outputs(4696) <= layer2_outputs(342);
    outputs(4697) <= not(layer2_outputs(3625));
    outputs(4698) <= layer2_outputs(2908);
    outputs(4699) <= not((layer2_outputs(8271)) and (layer2_outputs(7661)));
    outputs(4700) <= layer2_outputs(6667);
    outputs(4701) <= not(layer2_outputs(4469));
    outputs(4702) <= (layer2_outputs(1295)) and not (layer2_outputs(5708));
    outputs(4703) <= layer2_outputs(9913);
    outputs(4704) <= not(layer2_outputs(7426)) or (layer2_outputs(7651));
    outputs(4705) <= not((layer2_outputs(5050)) or (layer2_outputs(8551)));
    outputs(4706) <= (layer2_outputs(3505)) and (layer2_outputs(10122));
    outputs(4707) <= not(layer2_outputs(1169));
    outputs(4708) <= not(layer2_outputs(7664));
    outputs(4709) <= not(layer2_outputs(2400));
    outputs(4710) <= (layer2_outputs(7771)) xor (layer2_outputs(7906));
    outputs(4711) <= not(layer2_outputs(7204));
    outputs(4712) <= not(layer2_outputs(8823));
    outputs(4713) <= not(layer2_outputs(203));
    outputs(4714) <= layer2_outputs(3892);
    outputs(4715) <= layer2_outputs(3724);
    outputs(4716) <= not((layer2_outputs(8859)) xor (layer2_outputs(8042)));
    outputs(4717) <= layer2_outputs(9863);
    outputs(4718) <= (layer2_outputs(8827)) and not (layer2_outputs(7299));
    outputs(4719) <= (layer2_outputs(625)) and (layer2_outputs(7098));
    outputs(4720) <= not(layer2_outputs(4001)) or (layer2_outputs(409));
    outputs(4721) <= not(layer2_outputs(3641));
    outputs(4722) <= layer2_outputs(1969);
    outputs(4723) <= (layer2_outputs(3342)) and (layer2_outputs(5392));
    outputs(4724) <= not(layer2_outputs(2271));
    outputs(4725) <= layer2_outputs(4422);
    outputs(4726) <= not(layer2_outputs(8517));
    outputs(4727) <= not((layer2_outputs(63)) xor (layer2_outputs(2781)));
    outputs(4728) <= layer2_outputs(9790);
    outputs(4729) <= not((layer2_outputs(8566)) and (layer2_outputs(5593)));
    outputs(4730) <= layer2_outputs(9902);
    outputs(4731) <= not((layer2_outputs(975)) xor (layer2_outputs(9015)));
    outputs(4732) <= not(layer2_outputs(293));
    outputs(4733) <= layer2_outputs(4767);
    outputs(4734) <= (layer2_outputs(5718)) xor (layer2_outputs(5132));
    outputs(4735) <= not(layer2_outputs(1995)) or (layer2_outputs(9541));
    outputs(4736) <= not(layer2_outputs(7010));
    outputs(4737) <= not(layer2_outputs(9274));
    outputs(4738) <= not(layer2_outputs(2639));
    outputs(4739) <= (layer2_outputs(2537)) xor (layer2_outputs(5619));
    outputs(4740) <= not((layer2_outputs(9423)) xor (layer2_outputs(4655)));
    outputs(4741) <= (layer2_outputs(5544)) xor (layer2_outputs(1203));
    outputs(4742) <= (layer2_outputs(2647)) and not (layer2_outputs(1707));
    outputs(4743) <= layer2_outputs(8562);
    outputs(4744) <= layer2_outputs(3257);
    outputs(4745) <= not((layer2_outputs(6524)) xor (layer2_outputs(4657)));
    outputs(4746) <= (layer2_outputs(65)) or (layer2_outputs(8548));
    outputs(4747) <= not((layer2_outputs(8444)) xor (layer2_outputs(8866)));
    outputs(4748) <= not(layer2_outputs(6013));
    outputs(4749) <= (layer2_outputs(8567)) xor (layer2_outputs(2886));
    outputs(4750) <= (layer2_outputs(6563)) and (layer2_outputs(3857));
    outputs(4751) <= (layer2_outputs(1757)) xor (layer2_outputs(2370));
    outputs(4752) <= not(layer2_outputs(119));
    outputs(4753) <= not((layer2_outputs(1798)) xor (layer2_outputs(3494)));
    outputs(4754) <= not((layer2_outputs(5512)) xor (layer2_outputs(4613)));
    outputs(4755) <= layer2_outputs(5578);
    outputs(4756) <= not(layer2_outputs(6765));
    outputs(4757) <= layer2_outputs(91);
    outputs(4758) <= layer2_outputs(5631);
    outputs(4759) <= not(layer2_outputs(8598));
    outputs(4760) <= not((layer2_outputs(4473)) xor (layer2_outputs(9595)));
    outputs(4761) <= layer2_outputs(1465);
    outputs(4762) <= not((layer2_outputs(4760)) xor (layer2_outputs(6695)));
    outputs(4763) <= layer2_outputs(2775);
    outputs(4764) <= (layer2_outputs(2853)) xor (layer2_outputs(8013));
    outputs(4765) <= layer2_outputs(7827);
    outputs(4766) <= not(layer2_outputs(4824)) or (layer2_outputs(6157));
    outputs(4767) <= (layer2_outputs(3514)) and (layer2_outputs(6495));
    outputs(4768) <= not((layer2_outputs(9285)) xor (layer2_outputs(5525)));
    outputs(4769) <= (layer2_outputs(5221)) xor (layer2_outputs(9935));
    outputs(4770) <= not(layer2_outputs(4566));
    outputs(4771) <= (layer2_outputs(6866)) xor (layer2_outputs(2686));
    outputs(4772) <= (layer2_outputs(2075)) and (layer2_outputs(8716));
    outputs(4773) <= (layer2_outputs(420)) xor (layer2_outputs(7258));
    outputs(4774) <= layer2_outputs(7569);
    outputs(4775) <= not(layer2_outputs(8320));
    outputs(4776) <= layer2_outputs(8351);
    outputs(4777) <= layer2_outputs(3490);
    outputs(4778) <= (layer2_outputs(3684)) and (layer2_outputs(2605));
    outputs(4779) <= not((layer2_outputs(8711)) xor (layer2_outputs(8076)));
    outputs(4780) <= layer2_outputs(7180);
    outputs(4781) <= not(layer2_outputs(5520));
    outputs(4782) <= not((layer2_outputs(3939)) or (layer2_outputs(9153)));
    outputs(4783) <= layer2_outputs(4407);
    outputs(4784) <= not(layer2_outputs(5787));
    outputs(4785) <= layer2_outputs(3771);
    outputs(4786) <= layer2_outputs(1265);
    outputs(4787) <= (layer2_outputs(470)) and not (layer2_outputs(10238));
    outputs(4788) <= layer2_outputs(6550);
    outputs(4789) <= not((layer2_outputs(5957)) or (layer2_outputs(3157)));
    outputs(4790) <= not((layer2_outputs(3038)) xor (layer2_outputs(7321)));
    outputs(4791) <= layer2_outputs(4802);
    outputs(4792) <= (layer2_outputs(4343)) and not (layer2_outputs(5432));
    outputs(4793) <= (layer2_outputs(4808)) or (layer2_outputs(7320));
    outputs(4794) <= not(layer2_outputs(4547));
    outputs(4795) <= not((layer2_outputs(4095)) xor (layer2_outputs(6575)));
    outputs(4796) <= not(layer2_outputs(9669));
    outputs(4797) <= (layer2_outputs(2312)) xor (layer2_outputs(10185));
    outputs(4798) <= layer2_outputs(7759);
    outputs(4799) <= not(layer2_outputs(4355)) or (layer2_outputs(7008));
    outputs(4800) <= not((layer2_outputs(5398)) or (layer2_outputs(9811)));
    outputs(4801) <= layer2_outputs(7563);
    outputs(4802) <= not((layer2_outputs(7333)) or (layer2_outputs(5029)));
    outputs(4803) <= not(layer2_outputs(8780));
    outputs(4804) <= not(layer2_outputs(749));
    outputs(4805) <= not(layer2_outputs(8172));
    outputs(4806) <= not(layer2_outputs(4974));
    outputs(4807) <= not(layer2_outputs(3801));
    outputs(4808) <= not(layer2_outputs(9527)) or (layer2_outputs(6914));
    outputs(4809) <= (layer2_outputs(6922)) or (layer2_outputs(1355));
    outputs(4810) <= not((layer2_outputs(1803)) and (layer2_outputs(812)));
    outputs(4811) <= not(layer2_outputs(3531));
    outputs(4812) <= not((layer2_outputs(5078)) xor (layer2_outputs(1499)));
    outputs(4813) <= not((layer2_outputs(4655)) xor (layer2_outputs(4185)));
    outputs(4814) <= layer2_outputs(8020);
    outputs(4815) <= not(layer2_outputs(7662)) or (layer2_outputs(5638));
    outputs(4816) <= layer2_outputs(5515);
    outputs(4817) <= not((layer2_outputs(7930)) xor (layer2_outputs(2831)));
    outputs(4818) <= not(layer2_outputs(2531));
    outputs(4819) <= (layer2_outputs(8926)) and not (layer2_outputs(2623));
    outputs(4820) <= layer2_outputs(7493);
    outputs(4821) <= (layer2_outputs(35)) and (layer2_outputs(3747));
    outputs(4822) <= not(layer2_outputs(5447));
    outputs(4823) <= not(layer2_outputs(9547));
    outputs(4824) <= not(layer2_outputs(4724));
    outputs(4825) <= layer2_outputs(6622);
    outputs(4826) <= layer2_outputs(8276);
    outputs(4827) <= layer2_outputs(5812);
    outputs(4828) <= not(layer2_outputs(4880));
    outputs(4829) <= not((layer2_outputs(197)) or (layer2_outputs(7994)));
    outputs(4830) <= not(layer2_outputs(80));
    outputs(4831) <= layer2_outputs(9954);
    outputs(4832) <= not(layer2_outputs(8890));
    outputs(4833) <= not(layer2_outputs(8323));
    outputs(4834) <= (layer2_outputs(9613)) and not (layer2_outputs(1662));
    outputs(4835) <= not(layer2_outputs(8921));
    outputs(4836) <= not(layer2_outputs(3232));
    outputs(4837) <= layer2_outputs(7933);
    outputs(4838) <= not((layer2_outputs(694)) and (layer2_outputs(9084)));
    outputs(4839) <= not((layer2_outputs(1310)) or (layer2_outputs(18)));
    outputs(4840) <= layer2_outputs(4461);
    outputs(4841) <= not(layer2_outputs(665));
    outputs(4842) <= not(layer2_outputs(6735));
    outputs(4843) <= not((layer2_outputs(2293)) xor (layer2_outputs(4049)));
    outputs(4844) <= layer2_outputs(2968);
    outputs(4845) <= not(layer2_outputs(7013));
    outputs(4846) <= layer2_outputs(4107);
    outputs(4847) <= layer2_outputs(9853);
    outputs(4848) <= (layer2_outputs(4102)) and not (layer2_outputs(3241));
    outputs(4849) <= not((layer2_outputs(2803)) xor (layer2_outputs(1665)));
    outputs(4850) <= not(layer2_outputs(10169));
    outputs(4851) <= (layer2_outputs(7348)) and not (layer2_outputs(1599));
    outputs(4852) <= (layer2_outputs(9920)) and not (layer2_outputs(8033));
    outputs(4853) <= not((layer2_outputs(5151)) xor (layer2_outputs(4803)));
    outputs(4854) <= not((layer2_outputs(991)) xor (layer2_outputs(7271)));
    outputs(4855) <= (layer2_outputs(9863)) and not (layer2_outputs(3579));
    outputs(4856) <= not(layer2_outputs(9340)) or (layer2_outputs(1867));
    outputs(4857) <= not((layer2_outputs(3902)) xor (layer2_outputs(1991)));
    outputs(4858) <= not(layer2_outputs(1411));
    outputs(4859) <= not(layer2_outputs(4490));
    outputs(4860) <= not(layer2_outputs(9238)) or (layer2_outputs(613));
    outputs(4861) <= not(layer2_outputs(6486));
    outputs(4862) <= layer2_outputs(5144);
    outputs(4863) <= not(layer2_outputs(6740));
    outputs(4864) <= not((layer2_outputs(4734)) xor (layer2_outputs(8591)));
    outputs(4865) <= (layer2_outputs(5455)) xor (layer2_outputs(2401));
    outputs(4866) <= layer2_outputs(6426);
    outputs(4867) <= layer2_outputs(1987);
    outputs(4868) <= layer2_outputs(8564);
    outputs(4869) <= not((layer2_outputs(208)) xor (layer2_outputs(3808)));
    outputs(4870) <= (layer2_outputs(6995)) xor (layer2_outputs(5446));
    outputs(4871) <= not(layer2_outputs(9755));
    outputs(4872) <= (layer2_outputs(4136)) and not (layer2_outputs(5689));
    outputs(4873) <= layer2_outputs(9133);
    outputs(4874) <= not(layer2_outputs(737));
    outputs(4875) <= (layer2_outputs(4523)) and (layer2_outputs(568));
    outputs(4876) <= layer2_outputs(7112);
    outputs(4877) <= layer2_outputs(2912);
    outputs(4878) <= not(layer2_outputs(8782));
    outputs(4879) <= layer2_outputs(9731);
    outputs(4880) <= not((layer2_outputs(4913)) xor (layer2_outputs(9971)));
    outputs(4881) <= not((layer2_outputs(9390)) xor (layer2_outputs(7614)));
    outputs(4882) <= not(layer2_outputs(9051)) or (layer2_outputs(897));
    outputs(4883) <= (layer2_outputs(8337)) xor (layer2_outputs(5872));
    outputs(4884) <= not(layer2_outputs(4744));
    outputs(4885) <= not(layer2_outputs(2553));
    outputs(4886) <= (layer2_outputs(3379)) xor (layer2_outputs(1424));
    outputs(4887) <= (layer2_outputs(193)) xor (layer2_outputs(8273));
    outputs(4888) <= not(layer2_outputs(8026)) or (layer2_outputs(7103));
    outputs(4889) <= (layer2_outputs(4153)) or (layer2_outputs(2002));
    outputs(4890) <= (layer2_outputs(989)) xor (layer2_outputs(2783));
    outputs(4891) <= layer2_outputs(5102);
    outputs(4892) <= layer2_outputs(1796);
    outputs(4893) <= not(layer2_outputs(10095)) or (layer2_outputs(10007));
    outputs(4894) <= (layer2_outputs(10054)) xor (layer2_outputs(2275));
    outputs(4895) <= (layer2_outputs(4394)) xor (layer2_outputs(5489));
    outputs(4896) <= not(layer2_outputs(8990)) or (layer2_outputs(2311));
    outputs(4897) <= layer2_outputs(4607);
    outputs(4898) <= (layer2_outputs(10221)) and not (layer2_outputs(2375));
    outputs(4899) <= (layer2_outputs(2017)) and not (layer2_outputs(1207));
    outputs(4900) <= not(layer2_outputs(4761));
    outputs(4901) <= (layer2_outputs(9124)) and (layer2_outputs(2937));
    outputs(4902) <= not(layer2_outputs(8528));
    outputs(4903) <= (layer2_outputs(849)) and not (layer2_outputs(1522));
    outputs(4904) <= layer2_outputs(5462);
    outputs(4905) <= layer2_outputs(2748);
    outputs(4906) <= layer2_outputs(9961);
    outputs(4907) <= (layer2_outputs(5110)) xor (layer2_outputs(9753));
    outputs(4908) <= not(layer2_outputs(677));
    outputs(4909) <= not((layer2_outputs(6047)) xor (layer2_outputs(9176)));
    outputs(4910) <= not(layer2_outputs(640));
    outputs(4911) <= layer2_outputs(6019);
    outputs(4912) <= layer2_outputs(6316);
    outputs(4913) <= not(layer2_outputs(8144));
    outputs(4914) <= (layer2_outputs(622)) and not (layer2_outputs(3119));
    outputs(4915) <= layer2_outputs(5421);
    outputs(4916) <= layer2_outputs(2523);
    outputs(4917) <= not(layer2_outputs(2047));
    outputs(4918) <= layer2_outputs(2103);
    outputs(4919) <= not(layer2_outputs(7498));
    outputs(4920) <= not((layer2_outputs(884)) xor (layer2_outputs(2441)));
    outputs(4921) <= layer2_outputs(3841);
    outputs(4922) <= not(layer2_outputs(602));
    outputs(4923) <= (layer2_outputs(9918)) xor (layer2_outputs(1864));
    outputs(4924) <= not(layer2_outputs(314));
    outputs(4925) <= layer2_outputs(2625);
    outputs(4926) <= not(layer2_outputs(2372));
    outputs(4927) <= layer2_outputs(3782);
    outputs(4928) <= (layer2_outputs(5019)) and not (layer2_outputs(3732));
    outputs(4929) <= (layer2_outputs(7486)) and not (layer2_outputs(267));
    outputs(4930) <= layer2_outputs(3959);
    outputs(4931) <= (layer2_outputs(1489)) and (layer2_outputs(5431));
    outputs(4932) <= not((layer2_outputs(7329)) xor (layer2_outputs(9879)));
    outputs(4933) <= not(layer2_outputs(2443));
    outputs(4934) <= not(layer2_outputs(7652));
    outputs(4935) <= layer2_outputs(9533);
    outputs(4936) <= layer2_outputs(1659);
    outputs(4937) <= not(layer2_outputs(8664)) or (layer2_outputs(7900));
    outputs(4938) <= not(layer2_outputs(3538)) or (layer2_outputs(8177));
    outputs(4939) <= not(layer2_outputs(8530));
    outputs(4940) <= (layer2_outputs(5199)) and not (layer2_outputs(995));
    outputs(4941) <= not((layer2_outputs(5184)) or (layer2_outputs(8509)));
    outputs(4942) <= not((layer2_outputs(4290)) and (layer2_outputs(1215)));
    outputs(4943) <= not((layer2_outputs(8640)) or (layer2_outputs(7632)));
    outputs(4944) <= not(layer2_outputs(6367));
    outputs(4945) <= not((layer2_outputs(9875)) or (layer2_outputs(972)));
    outputs(4946) <= not(layer2_outputs(7368));
    outputs(4947) <= not(layer2_outputs(3331));
    outputs(4948) <= (layer2_outputs(7271)) and not (layer2_outputs(739));
    outputs(4949) <= (layer2_outputs(8558)) and not (layer2_outputs(5327));
    outputs(4950) <= not(layer2_outputs(6021));
    outputs(4951) <= (layer2_outputs(6469)) or (layer2_outputs(3411));
    outputs(4952) <= layer2_outputs(623);
    outputs(4953) <= (layer2_outputs(1816)) and (layer2_outputs(6734));
    outputs(4954) <= (layer2_outputs(2382)) and (layer2_outputs(4955));
    outputs(4955) <= not((layer2_outputs(6527)) or (layer2_outputs(0)));
    outputs(4956) <= (layer2_outputs(1405)) xor (layer2_outputs(3376));
    outputs(4957) <= not(layer2_outputs(8836));
    outputs(4958) <= not(layer2_outputs(1541));
    outputs(4959) <= not(layer2_outputs(7525)) or (layer2_outputs(6395));
    outputs(4960) <= not(layer2_outputs(8670));
    outputs(4961) <= (layer2_outputs(5480)) xor (layer2_outputs(3056));
    outputs(4962) <= (layer2_outputs(9800)) and not (layer2_outputs(5051));
    outputs(4963) <= (layer2_outputs(3619)) or (layer2_outputs(9696));
    outputs(4964) <= layer2_outputs(2391);
    outputs(4965) <= not(layer2_outputs(7709));
    outputs(4966) <= layer2_outputs(7219);
    outputs(4967) <= layer2_outputs(9432);
    outputs(4968) <= layer2_outputs(7017);
    outputs(4969) <= not((layer2_outputs(2705)) and (layer2_outputs(5934)));
    outputs(4970) <= not(layer2_outputs(3983));
    outputs(4971) <= layer2_outputs(8461);
    outputs(4972) <= (layer2_outputs(5648)) and not (layer2_outputs(2671));
    outputs(4973) <= not(layer2_outputs(9430));
    outputs(4974) <= (layer2_outputs(2729)) xor (layer2_outputs(763));
    outputs(4975) <= not(layer2_outputs(1439));
    outputs(4976) <= not((layer2_outputs(2713)) or (layer2_outputs(7667)));
    outputs(4977) <= not(layer2_outputs(922));
    outputs(4978) <= layer2_outputs(3207);
    outputs(4979) <= not((layer2_outputs(3767)) or (layer2_outputs(3915)));
    outputs(4980) <= not(layer2_outputs(4963));
    outputs(4981) <= (layer2_outputs(4295)) and not (layer2_outputs(2420));
    outputs(4982) <= not((layer2_outputs(662)) xor (layer2_outputs(6757)));
    outputs(4983) <= layer2_outputs(930);
    outputs(4984) <= not((layer2_outputs(1909)) xor (layer2_outputs(9880)));
    outputs(4985) <= layer2_outputs(9786);
    outputs(4986) <= (layer2_outputs(4181)) xor (layer2_outputs(1082));
    outputs(4987) <= layer2_outputs(7659);
    outputs(4988) <= not(layer2_outputs(10044));
    outputs(4989) <= not(layer2_outputs(5755));
    outputs(4990) <= not(layer2_outputs(5419)) or (layer2_outputs(5764));
    outputs(4991) <= layer2_outputs(8071);
    outputs(4992) <= not(layer2_outputs(4695));
    outputs(4993) <= not(layer2_outputs(3367)) or (layer2_outputs(10168));
    outputs(4994) <= not(layer2_outputs(5275)) or (layer2_outputs(8802));
    outputs(4995) <= not(layer2_outputs(1518));
    outputs(4996) <= not(layer2_outputs(5546)) or (layer2_outputs(809));
    outputs(4997) <= not(layer2_outputs(6466));
    outputs(4998) <= (layer2_outputs(9172)) xor (layer2_outputs(924));
    outputs(4999) <= not((layer2_outputs(7689)) xor (layer2_outputs(30)));
    outputs(5000) <= layer2_outputs(140);
    outputs(5001) <= not(layer2_outputs(4745));
    outputs(5002) <= not((layer2_outputs(6118)) xor (layer2_outputs(7528)));
    outputs(5003) <= not((layer2_outputs(3758)) xor (layer2_outputs(2421)));
    outputs(5004) <= layer2_outputs(3835);
    outputs(5005) <= not(layer2_outputs(8408));
    outputs(5006) <= not(layer2_outputs(9635));
    outputs(5007) <= not(layer2_outputs(2549));
    outputs(5008) <= layer2_outputs(3360);
    outputs(5009) <= (layer2_outputs(2711)) xor (layer2_outputs(6156));
    outputs(5010) <= not(layer2_outputs(5810));
    outputs(5011) <= (layer2_outputs(7369)) and not (layer2_outputs(3568));
    outputs(5012) <= (layer2_outputs(8394)) xor (layer2_outputs(8891));
    outputs(5013) <= layer2_outputs(2831);
    outputs(5014) <= not(layer2_outputs(2040));
    outputs(5015) <= (layer2_outputs(5877)) and (layer2_outputs(10018));
    outputs(5016) <= not(layer2_outputs(5581)) or (layer2_outputs(5878));
    outputs(5017) <= not((layer2_outputs(5820)) or (layer2_outputs(5052)));
    outputs(5018) <= not(layer2_outputs(8761)) or (layer2_outputs(5033));
    outputs(5019) <= layer2_outputs(5950);
    outputs(5020) <= not(layer2_outputs(9839));
    outputs(5021) <= layer2_outputs(5307);
    outputs(5022) <= not((layer2_outputs(3353)) and (layer2_outputs(8524)));
    outputs(5023) <= not(layer2_outputs(4909));
    outputs(5024) <= (layer2_outputs(4824)) xor (layer2_outputs(5669));
    outputs(5025) <= layer2_outputs(5256);
    outputs(5026) <= not(layer2_outputs(3927));
    outputs(5027) <= layer2_outputs(2505);
    outputs(5028) <= not(layer2_outputs(8610));
    outputs(5029) <= layer2_outputs(3958);
    outputs(5030) <= layer2_outputs(9441);
    outputs(5031) <= not(layer2_outputs(4111));
    outputs(5032) <= not((layer2_outputs(7060)) and (layer2_outputs(1749)));
    outputs(5033) <= not(layer2_outputs(6216)) or (layer2_outputs(1243));
    outputs(5034) <= (layer2_outputs(7082)) and not (layer2_outputs(6913));
    outputs(5035) <= not(layer2_outputs(10012)) or (layer2_outputs(6689));
    outputs(5036) <= (layer2_outputs(10019)) xor (layer2_outputs(1997));
    outputs(5037) <= not(layer2_outputs(1018));
    outputs(5038) <= not(layer2_outputs(344)) or (layer2_outputs(2899));
    outputs(5039) <= not(layer2_outputs(3844));
    outputs(5040) <= (layer2_outputs(4335)) and not (layer2_outputs(1273));
    outputs(5041) <= (layer2_outputs(9265)) and not (layer2_outputs(2557));
    outputs(5042) <= not(layer2_outputs(2905));
    outputs(5043) <= layer2_outputs(9463);
    outputs(5044) <= not((layer2_outputs(7551)) or (layer2_outputs(979)));
    outputs(5045) <= layer2_outputs(7261);
    outputs(5046) <= (layer2_outputs(4658)) and (layer2_outputs(5040));
    outputs(5047) <= layer2_outputs(3220);
    outputs(5048) <= (layer2_outputs(4190)) xor (layer2_outputs(4003));
    outputs(5049) <= not(layer2_outputs(5545));
    outputs(5050) <= not((layer2_outputs(10064)) xor (layer2_outputs(825)));
    outputs(5051) <= layer2_outputs(8194);
    outputs(5052) <= layer2_outputs(5197);
    outputs(5053) <= not(layer2_outputs(1344));
    outputs(5054) <= not(layer2_outputs(523));
    outputs(5055) <= not(layer2_outputs(920));
    outputs(5056) <= not((layer2_outputs(6002)) xor (layer2_outputs(562)));
    outputs(5057) <= not(layer2_outputs(7627));
    outputs(5058) <= layer2_outputs(8232);
    outputs(5059) <= not(layer2_outputs(8789));
    outputs(5060) <= not(layer2_outputs(8850));
    outputs(5061) <= layer2_outputs(3843);
    outputs(5062) <= not(layer2_outputs(8829));
    outputs(5063) <= not(layer2_outputs(10059)) or (layer2_outputs(5965));
    outputs(5064) <= layer2_outputs(5561);
    outputs(5065) <= not(layer2_outputs(7056));
    outputs(5066) <= layer2_outputs(1619);
    outputs(5067) <= not(layer2_outputs(5081));
    outputs(5068) <= not((layer2_outputs(5936)) xor (layer2_outputs(6787)));
    outputs(5069) <= not((layer2_outputs(1177)) or (layer2_outputs(7951)));
    outputs(5070) <= (layer2_outputs(7904)) and (layer2_outputs(93));
    outputs(5071) <= (layer2_outputs(4879)) xor (layer2_outputs(10213));
    outputs(5072) <= not(layer2_outputs(5315));
    outputs(5073) <= (layer2_outputs(9557)) xor (layer2_outputs(1859));
    outputs(5074) <= (layer2_outputs(5933)) xor (layer2_outputs(9016));
    outputs(5075) <= (layer2_outputs(4445)) xor (layer2_outputs(3965));
    outputs(5076) <= not((layer2_outputs(5700)) xor (layer2_outputs(9651)));
    outputs(5077) <= not((layer2_outputs(2612)) or (layer2_outputs(5100)));
    outputs(5078) <= (layer2_outputs(2625)) xor (layer2_outputs(7860));
    outputs(5079) <= not(layer2_outputs(5203)) or (layer2_outputs(5925));
    outputs(5080) <= not(layer2_outputs(6837));
    outputs(5081) <= layer2_outputs(2763);
    outputs(5082) <= not(layer2_outputs(5189));
    outputs(5083) <= not(layer2_outputs(10187));
    outputs(5084) <= not((layer2_outputs(8109)) xor (layer2_outputs(6677)));
    outputs(5085) <= not(layer2_outputs(6844));
    outputs(5086) <= layer2_outputs(8192);
    outputs(5087) <= layer2_outputs(8013);
    outputs(5088) <= not(layer2_outputs(9049)) or (layer2_outputs(1325));
    outputs(5089) <= not(layer2_outputs(903));
    outputs(5090) <= not(layer2_outputs(2867));
    outputs(5091) <= not(layer2_outputs(7672));
    outputs(5092) <= layer2_outputs(1157);
    outputs(5093) <= layer2_outputs(5902);
    outputs(5094) <= layer2_outputs(6841);
    outputs(5095) <= (layer2_outputs(5881)) or (layer2_outputs(1601));
    outputs(5096) <= not(layer2_outputs(3426));
    outputs(5097) <= not(layer2_outputs(5794));
    outputs(5098) <= not((layer2_outputs(6364)) or (layer2_outputs(4367)));
    outputs(5099) <= not(layer2_outputs(9130)) or (layer2_outputs(1892));
    outputs(5100) <= not(layer2_outputs(9508));
    outputs(5101) <= layer2_outputs(3123);
    outputs(5102) <= layer2_outputs(2085);
    outputs(5103) <= (layer2_outputs(1346)) and not (layer2_outputs(9204));
    outputs(5104) <= not((layer2_outputs(2529)) xor (layer2_outputs(6098)));
    outputs(5105) <= not(layer2_outputs(1637)) or (layer2_outputs(1303));
    outputs(5106) <= (layer2_outputs(9090)) xor (layer2_outputs(2265));
    outputs(5107) <= layer2_outputs(7127);
    outputs(5108) <= not((layer2_outputs(2767)) xor (layer2_outputs(5182)));
    outputs(5109) <= not(layer2_outputs(799)) or (layer2_outputs(780));
    outputs(5110) <= layer2_outputs(7520);
    outputs(5111) <= (layer2_outputs(7819)) xor (layer2_outputs(7081));
    outputs(5112) <= not(layer2_outputs(5632));
    outputs(5113) <= not(layer2_outputs(9751));
    outputs(5114) <= not(layer2_outputs(6796));
    outputs(5115) <= not((layer2_outputs(6033)) or (layer2_outputs(1421)));
    outputs(5116) <= (layer2_outputs(6709)) and (layer2_outputs(3452));
    outputs(5117) <= layer2_outputs(5654);
    outputs(5118) <= not(layer2_outputs(1506));
    outputs(5119) <= not(layer2_outputs(3991));
    outputs(5120) <= not(layer2_outputs(6299));
    outputs(5121) <= not(layer2_outputs(4250)) or (layer2_outputs(1755));
    outputs(5122) <= (layer2_outputs(9568)) xor (layer2_outputs(9475));
    outputs(5123) <= not((layer2_outputs(3179)) xor (layer2_outputs(4240)));
    outputs(5124) <= not(layer2_outputs(9877));
    outputs(5125) <= (layer2_outputs(2462)) and not (layer2_outputs(8901));
    outputs(5126) <= layer2_outputs(9448);
    outputs(5127) <= (layer2_outputs(1737)) xor (layer2_outputs(2207));
    outputs(5128) <= not((layer2_outputs(6029)) xor (layer2_outputs(2860)));
    outputs(5129) <= (layer2_outputs(9949)) xor (layer2_outputs(4607));
    outputs(5130) <= (layer2_outputs(4042)) xor (layer2_outputs(6357));
    outputs(5131) <= layer2_outputs(8652);
    outputs(5132) <= layer2_outputs(1628);
    outputs(5133) <= layer2_outputs(3697);
    outputs(5134) <= not(layer2_outputs(668));
    outputs(5135) <= not(layer2_outputs(3345));
    outputs(5136) <= not(layer2_outputs(8215));
    outputs(5137) <= not((layer2_outputs(5670)) xor (layer2_outputs(10182)));
    outputs(5138) <= (layer2_outputs(5408)) or (layer2_outputs(3335));
    outputs(5139) <= not(layer2_outputs(1052));
    outputs(5140) <= not((layer2_outputs(6079)) xor (layer2_outputs(10234)));
    outputs(5141) <= (layer2_outputs(4365)) xor (layer2_outputs(541));
    outputs(5142) <= layer2_outputs(5786);
    outputs(5143) <= not(layer2_outputs(9417)) or (layer2_outputs(47));
    outputs(5144) <= not(layer2_outputs(8561));
    outputs(5145) <= layer2_outputs(6169);
    outputs(5146) <= not(layer2_outputs(9666)) or (layer2_outputs(703));
    outputs(5147) <= not((layer2_outputs(7794)) xor (layer2_outputs(2528)));
    outputs(5148) <= (layer2_outputs(7767)) xor (layer2_outputs(9154));
    outputs(5149) <= (layer2_outputs(3435)) and (layer2_outputs(819));
    outputs(5150) <= (layer2_outputs(6547)) and not (layer2_outputs(8900));
    outputs(5151) <= not((layer2_outputs(268)) xor (layer2_outputs(5104)));
    outputs(5152) <= not((layer2_outputs(2639)) xor (layer2_outputs(5414)));
    outputs(5153) <= layer2_outputs(3616);
    outputs(5154) <= not(layer2_outputs(6844));
    outputs(5155) <= layer2_outputs(5030);
    outputs(5156) <= (layer2_outputs(8809)) or (layer2_outputs(9532));
    outputs(5157) <= (layer2_outputs(10206)) xor (layer2_outputs(3612));
    outputs(5158) <= not(layer2_outputs(2689)) or (layer2_outputs(9302));
    outputs(5159) <= layer2_outputs(381);
    outputs(5160) <= not(layer2_outputs(1710));
    outputs(5161) <= not(layer2_outputs(9663));
    outputs(5162) <= not((layer2_outputs(6204)) xor (layer2_outputs(8861)));
    outputs(5163) <= (layer2_outputs(829)) and (layer2_outputs(6768));
    outputs(5164) <= layer2_outputs(9565);
    outputs(5165) <= (layer2_outputs(5180)) and (layer2_outputs(9063));
    outputs(5166) <= not(layer2_outputs(6028));
    outputs(5167) <= not(layer2_outputs(4920)) or (layer2_outputs(9497));
    outputs(5168) <= layer2_outputs(929);
    outputs(5169) <= not((layer2_outputs(7320)) xor (layer2_outputs(2621)));
    outputs(5170) <= not(layer2_outputs(9281));
    outputs(5171) <= (layer2_outputs(5040)) and not (layer2_outputs(6014));
    outputs(5172) <= not(layer2_outputs(6327));
    outputs(5173) <= not(layer2_outputs(8439));
    outputs(5174) <= (layer2_outputs(6265)) xor (layer2_outputs(9736));
    outputs(5175) <= not((layer2_outputs(7703)) xor (layer2_outputs(4398)));
    outputs(5176) <= not(layer2_outputs(6620));
    outputs(5177) <= layer2_outputs(27);
    outputs(5178) <= not(layer2_outputs(7581));
    outputs(5179) <= not(layer2_outputs(4776));
    outputs(5180) <= layer2_outputs(8371);
    outputs(5181) <= layer2_outputs(5613);
    outputs(5182) <= layer2_outputs(2397);
    outputs(5183) <= not(layer2_outputs(7502));
    outputs(5184) <= not(layer2_outputs(9505));
    outputs(5185) <= not(layer2_outputs(7569));
    outputs(5186) <= not(layer2_outputs(2262));
    outputs(5187) <= layer2_outputs(20);
    outputs(5188) <= not((layer2_outputs(7377)) and (layer2_outputs(5502)));
    outputs(5189) <= not(layer2_outputs(4965));
    outputs(5190) <= (layer2_outputs(217)) xor (layer2_outputs(10166));
    outputs(5191) <= not(layer2_outputs(3464));
    outputs(5192) <= layer2_outputs(7323);
    outputs(5193) <= not(layer2_outputs(8858));
    outputs(5194) <= layer2_outputs(1324);
    outputs(5195) <= not(layer2_outputs(4910));
    outputs(5196) <= not(layer2_outputs(7869));
    outputs(5197) <= (layer2_outputs(7989)) xor (layer2_outputs(6043));
    outputs(5198) <= layer2_outputs(3320);
    outputs(5199) <= not(layer2_outputs(8425)) or (layer2_outputs(8002));
    outputs(5200) <= not(layer2_outputs(2375));
    outputs(5201) <= not(layer2_outputs(5537));
    outputs(5202) <= not(layer2_outputs(6237));
    outputs(5203) <= (layer2_outputs(7532)) xor (layer2_outputs(5099));
    outputs(5204) <= layer2_outputs(1861);
    outputs(5205) <= not(layer2_outputs(578));
    outputs(5206) <= not(layer2_outputs(7210));
    outputs(5207) <= not(layer2_outputs(2842));
    outputs(5208) <= not(layer2_outputs(2382));
    outputs(5209) <= not(layer2_outputs(8414));
    outputs(5210) <= not((layer2_outputs(3590)) xor (layer2_outputs(7934)));
    outputs(5211) <= not(layer2_outputs(7737));
    outputs(5212) <= layer2_outputs(6684);
    outputs(5213) <= not((layer2_outputs(2744)) xor (layer2_outputs(401)));
    outputs(5214) <= not((layer2_outputs(5516)) xor (layer2_outputs(6680)));
    outputs(5215) <= layer2_outputs(5829);
    outputs(5216) <= layer2_outputs(965);
    outputs(5217) <= not(layer2_outputs(1913));
    outputs(5218) <= (layer2_outputs(7822)) xor (layer2_outputs(6439));
    outputs(5219) <= layer2_outputs(6982);
    outputs(5220) <= not((layer2_outputs(1176)) xor (layer2_outputs(3388)));
    outputs(5221) <= not((layer2_outputs(1685)) xor (layer2_outputs(1633)));
    outputs(5222) <= (layer2_outputs(2233)) or (layer2_outputs(7766));
    outputs(5223) <= not((layer2_outputs(3288)) xor (layer2_outputs(3769)));
    outputs(5224) <= (layer2_outputs(9446)) xor (layer2_outputs(3195));
    outputs(5225) <= not(layer2_outputs(5226)) or (layer2_outputs(10132));
    outputs(5226) <= layer2_outputs(11);
    outputs(5227) <= layer2_outputs(9661);
    outputs(5228) <= not(layer2_outputs(7215));
    outputs(5229) <= (layer2_outputs(9360)) or (layer2_outputs(6083));
    outputs(5230) <= layer2_outputs(1533);
    outputs(5231) <= not((layer2_outputs(7090)) xor (layer2_outputs(9803)));
    outputs(5232) <= layer2_outputs(4504);
    outputs(5233) <= not(layer2_outputs(3381));
    outputs(5234) <= layer2_outputs(4828);
    outputs(5235) <= not((layer2_outputs(5370)) xor (layer2_outputs(2934)));
    outputs(5236) <= not((layer2_outputs(2187)) or (layer2_outputs(10195)));
    outputs(5237) <= layer2_outputs(1986);
    outputs(5238) <= (layer2_outputs(1628)) xor (layer2_outputs(5198));
    outputs(5239) <= layer2_outputs(6429);
    outputs(5240) <= not(layer2_outputs(1706)) or (layer2_outputs(6196));
    outputs(5241) <= layer2_outputs(7792);
    outputs(5242) <= not((layer2_outputs(620)) xor (layer2_outputs(8860)));
    outputs(5243) <= (layer2_outputs(7422)) xor (layer2_outputs(4661));
    outputs(5244) <= (layer2_outputs(5563)) xor (layer2_outputs(8025));
    outputs(5245) <= (layer2_outputs(9834)) and (layer2_outputs(965));
    outputs(5246) <= layer2_outputs(9494);
    outputs(5247) <= not(layer2_outputs(10116));
    outputs(5248) <= not((layer2_outputs(8235)) xor (layer2_outputs(9122)));
    outputs(5249) <= (layer2_outputs(1778)) and not (layer2_outputs(9495));
    outputs(5250) <= not(layer2_outputs(9208));
    outputs(5251) <= not(layer2_outputs(5566));
    outputs(5252) <= layer2_outputs(5109);
    outputs(5253) <= not(layer2_outputs(2545));
    outputs(5254) <= not((layer2_outputs(7424)) xor (layer2_outputs(3666)));
    outputs(5255) <= not(layer2_outputs(7591));
    outputs(5256) <= not(layer2_outputs(2598)) or (layer2_outputs(5982));
    outputs(5257) <= not((layer2_outputs(10175)) xor (layer2_outputs(4703)));
    outputs(5258) <= not((layer2_outputs(1385)) xor (layer2_outputs(2655)));
    outputs(5259) <= not(layer2_outputs(9775));
    outputs(5260) <= not(layer2_outputs(5148)) or (layer2_outputs(8532));
    outputs(5261) <= not((layer2_outputs(1493)) xor (layer2_outputs(8058)));
    outputs(5262) <= not(layer2_outputs(946));
    outputs(5263) <= not((layer2_outputs(6259)) or (layer2_outputs(7340)));
    outputs(5264) <= (layer2_outputs(1129)) xor (layer2_outputs(1938));
    outputs(5265) <= not((layer2_outputs(9998)) xor (layer2_outputs(8552)));
    outputs(5266) <= not(layer2_outputs(5069));
    outputs(5267) <= not((layer2_outputs(2326)) xor (layer2_outputs(3303)));
    outputs(5268) <= not(layer2_outputs(4506));
    outputs(5269) <= not((layer2_outputs(7282)) xor (layer2_outputs(8218)));
    outputs(5270) <= not(layer2_outputs(3993));
    outputs(5271) <= not(layer2_outputs(5884));
    outputs(5272) <= layer2_outputs(512);
    outputs(5273) <= layer2_outputs(4727);
    outputs(5274) <= layer2_outputs(6435);
    outputs(5275) <= (layer2_outputs(9719)) and not (layer2_outputs(6293));
    outputs(5276) <= (layer2_outputs(2943)) or (layer2_outputs(7447));
    outputs(5277) <= not(layer2_outputs(6850)) or (layer2_outputs(1487));
    outputs(5278) <= layer2_outputs(4535);
    outputs(5279) <= not(layer2_outputs(3011));
    outputs(5280) <= (layer2_outputs(4182)) and not (layer2_outputs(8526));
    outputs(5281) <= not(layer2_outputs(8909));
    outputs(5282) <= not(layer2_outputs(640));
    outputs(5283) <= (layer2_outputs(9239)) xor (layer2_outputs(3335));
    outputs(5284) <= not(layer2_outputs(1820));
    outputs(5285) <= (layer2_outputs(3947)) xor (layer2_outputs(4459));
    outputs(5286) <= layer2_outputs(7902);
    outputs(5287) <= not(layer2_outputs(4707));
    outputs(5288) <= layer2_outputs(457);
    outputs(5289) <= layer2_outputs(5695);
    outputs(5290) <= not((layer2_outputs(2422)) xor (layer2_outputs(9367)));
    outputs(5291) <= not((layer2_outputs(6593)) and (layer2_outputs(1953)));
    outputs(5292) <= not(layer2_outputs(8294));
    outputs(5293) <= (layer2_outputs(7981)) xor (layer2_outputs(8187));
    outputs(5294) <= (layer2_outputs(4636)) and not (layer2_outputs(22));
    outputs(5295) <= not((layer2_outputs(5738)) xor (layer2_outputs(6136)));
    outputs(5296) <= not(layer2_outputs(1460));
    outputs(5297) <= not(layer2_outputs(7594)) or (layer2_outputs(8051));
    outputs(5298) <= layer2_outputs(9628);
    outputs(5299) <= not(layer2_outputs(3034)) or (layer2_outputs(8413));
    outputs(5300) <= layer2_outputs(5092);
    outputs(5301) <= not(layer2_outputs(3290));
    outputs(5302) <= layer2_outputs(8832);
    outputs(5303) <= (layer2_outputs(7380)) and not (layer2_outputs(8226));
    outputs(5304) <= not(layer2_outputs(4317));
    outputs(5305) <= not(layer2_outputs(10061));
    outputs(5306) <= (layer2_outputs(6094)) and not (layer2_outputs(6974));
    outputs(5307) <= not(layer2_outputs(2714)) or (layer2_outputs(2702));
    outputs(5308) <= (layer2_outputs(6097)) xor (layer2_outputs(9617));
    outputs(5309) <= (layer2_outputs(4100)) and not (layer2_outputs(6880));
    outputs(5310) <= layer2_outputs(7311);
    outputs(5311) <= layer2_outputs(6076);
    outputs(5312) <= not(layer2_outputs(5813));
    outputs(5313) <= not((layer2_outputs(5108)) xor (layer2_outputs(7482)));
    outputs(5314) <= not(layer2_outputs(7591));
    outputs(5315) <= layer2_outputs(3308);
    outputs(5316) <= layer2_outputs(1184);
    outputs(5317) <= (layer2_outputs(1392)) or (layer2_outputs(8535));
    outputs(5318) <= (layer2_outputs(7837)) xor (layer2_outputs(9933));
    outputs(5319) <= layer2_outputs(5154);
    outputs(5320) <= (layer2_outputs(5291)) xor (layer2_outputs(5405));
    outputs(5321) <= not((layer2_outputs(5862)) xor (layer2_outputs(2936)));
    outputs(5322) <= layer2_outputs(6380);
    outputs(5323) <= (layer2_outputs(8327)) xor (layer2_outputs(4803));
    outputs(5324) <= layer2_outputs(2699);
    outputs(5325) <= not(layer2_outputs(1122));
    outputs(5326) <= not((layer2_outputs(8068)) xor (layer2_outputs(9587)));
    outputs(5327) <= (layer2_outputs(9447)) xor (layer2_outputs(9250));
    outputs(5328) <= (layer2_outputs(2914)) xor (layer2_outputs(7192));
    outputs(5329) <= not((layer2_outputs(236)) xor (layer2_outputs(8240)));
    outputs(5330) <= layer2_outputs(9998);
    outputs(5331) <= not(layer2_outputs(10139)) or (layer2_outputs(7784));
    outputs(5332) <= layer2_outputs(9342);
    outputs(5333) <= layer2_outputs(872);
    outputs(5334) <= not(layer2_outputs(4730));
    outputs(5335) <= not((layer2_outputs(4914)) xor (layer2_outputs(1970)));
    outputs(5336) <= not(layer2_outputs(2579));
    outputs(5337) <= not(layer2_outputs(432));
    outputs(5338) <= layer2_outputs(9302);
    outputs(5339) <= not((layer2_outputs(1095)) xor (layer2_outputs(8793)));
    outputs(5340) <= not(layer2_outputs(5200)) or (layer2_outputs(1553));
    outputs(5341) <= not(layer2_outputs(1887)) or (layer2_outputs(9353));
    outputs(5342) <= (layer2_outputs(623)) xor (layer2_outputs(7440));
    outputs(5343) <= layer2_outputs(3085);
    outputs(5344) <= not(layer2_outputs(2320));
    outputs(5345) <= layer2_outputs(2967);
    outputs(5346) <= not(layer2_outputs(9959));
    outputs(5347) <= layer2_outputs(4382);
    outputs(5348) <= layer2_outputs(1180);
    outputs(5349) <= layer2_outputs(451);
    outputs(5350) <= not(layer2_outputs(6820));
    outputs(5351) <= layer2_outputs(5205);
    outputs(5352) <= not(layer2_outputs(8111));
    outputs(5353) <= layer2_outputs(567);
    outputs(5354) <= (layer2_outputs(8002)) and not (layer2_outputs(5455));
    outputs(5355) <= (layer2_outputs(5751)) xor (layer2_outputs(3261));
    outputs(5356) <= layer2_outputs(9230);
    outputs(5357) <= not(layer2_outputs(75));
    outputs(5358) <= layer2_outputs(2576);
    outputs(5359) <= not(layer2_outputs(7252)) or (layer2_outputs(5690));
    outputs(5360) <= (layer2_outputs(23)) and (layer2_outputs(5918));
    outputs(5361) <= not(layer2_outputs(8710));
    outputs(5362) <= layer2_outputs(517);
    outputs(5363) <= not(layer2_outputs(1236));
    outputs(5364) <= (layer2_outputs(7345)) xor (layer2_outputs(8283));
    outputs(5365) <= not(layer2_outputs(5300));
    outputs(5366) <= (layer2_outputs(8621)) xor (layer2_outputs(5032));
    outputs(5367) <= (layer2_outputs(3673)) xor (layer2_outputs(903));
    outputs(5368) <= layer2_outputs(2559);
    outputs(5369) <= not((layer2_outputs(454)) xor (layer2_outputs(7065)));
    outputs(5370) <= not(layer2_outputs(9394));
    outputs(5371) <= not(layer2_outputs(5254));
    outputs(5372) <= (layer2_outputs(5100)) xor (layer2_outputs(4434));
    outputs(5373) <= not(layer2_outputs(1261));
    outputs(5374) <= (layer2_outputs(6628)) xor (layer2_outputs(8466));
    outputs(5375) <= not((layer2_outputs(7112)) xor (layer2_outputs(4942)));
    outputs(5376) <= (layer2_outputs(8066)) or (layer2_outputs(421));
    outputs(5377) <= not((layer2_outputs(5055)) xor (layer2_outputs(1146)));
    outputs(5378) <= not(layer2_outputs(836)) or (layer2_outputs(5632));
    outputs(5379) <= not(layer2_outputs(4621));
    outputs(5380) <= layer2_outputs(5211);
    outputs(5381) <= not((layer2_outputs(947)) and (layer2_outputs(8987)));
    outputs(5382) <= not((layer2_outputs(5222)) and (layer2_outputs(2670)));
    outputs(5383) <= layer2_outputs(1585);
    outputs(5384) <= (layer2_outputs(8997)) xor (layer2_outputs(9914));
    outputs(5385) <= not(layer2_outputs(6771));
    outputs(5386) <= layer2_outputs(4984);
    outputs(5387) <= layer2_outputs(3806);
    outputs(5388) <= layer2_outputs(4072);
    outputs(5389) <= not(layer2_outputs(8924));
    outputs(5390) <= (layer2_outputs(3973)) or (layer2_outputs(955));
    outputs(5391) <= (layer2_outputs(9120)) xor (layer2_outputs(7001));
    outputs(5392) <= (layer2_outputs(209)) xor (layer2_outputs(5991));
    outputs(5393) <= layer2_outputs(1163);
    outputs(5394) <= not((layer2_outputs(3936)) xor (layer2_outputs(5844)));
    outputs(5395) <= layer2_outputs(4430);
    outputs(5396) <= layer2_outputs(77);
    outputs(5397) <= not(layer2_outputs(7436));
    outputs(5398) <= layer2_outputs(7823);
    outputs(5399) <= (layer2_outputs(1378)) xor (layer2_outputs(6302));
    outputs(5400) <= layer2_outputs(7825);
    outputs(5401) <= layer2_outputs(192);
    outputs(5402) <= (layer2_outputs(517)) and (layer2_outputs(4684));
    outputs(5403) <= not(layer2_outputs(1746));
    outputs(5404) <= not((layer2_outputs(5598)) xor (layer2_outputs(3276)));
    outputs(5405) <= not(layer2_outputs(6923));
    outputs(5406) <= (layer2_outputs(7179)) xor (layer2_outputs(2339));
    outputs(5407) <= layer2_outputs(390);
    outputs(5408) <= not(layer2_outputs(3505)) or (layer2_outputs(696));
    outputs(5409) <= (layer2_outputs(6208)) and not (layer2_outputs(1731));
    outputs(5410) <= (layer2_outputs(1844)) xor (layer2_outputs(9568));
    outputs(5411) <= (layer2_outputs(10154)) xor (layer2_outputs(10186));
    outputs(5412) <= not(layer2_outputs(4156));
    outputs(5413) <= not(layer2_outputs(8944));
    outputs(5414) <= layer2_outputs(4683);
    outputs(5415) <= layer2_outputs(1047);
    outputs(5416) <= (layer2_outputs(9203)) xor (layer2_outputs(514));
    outputs(5417) <= layer2_outputs(189);
    outputs(5418) <= layer2_outputs(3212);
    outputs(5419) <= not((layer2_outputs(7859)) xor (layer2_outputs(6792)));
    outputs(5420) <= not((layer2_outputs(9571)) xor (layer2_outputs(9805)));
    outputs(5421) <= not(layer2_outputs(6322)) or (layer2_outputs(3158));
    outputs(5422) <= (layer2_outputs(4205)) xor (layer2_outputs(9303));
    outputs(5423) <= (layer2_outputs(669)) and not (layer2_outputs(7742));
    outputs(5424) <= not(layer2_outputs(9495));
    outputs(5425) <= not(layer2_outputs(6341));
    outputs(5426) <= (layer2_outputs(59)) xor (layer2_outputs(3488));
    outputs(5427) <= layer2_outputs(92);
    outputs(5428) <= not(layer2_outputs(6906)) or (layer2_outputs(4654));
    outputs(5429) <= (layer2_outputs(5671)) xor (layer2_outputs(4083));
    outputs(5430) <= not((layer2_outputs(1498)) xor (layer2_outputs(5185)));
    outputs(5431) <= not((layer2_outputs(423)) xor (layer2_outputs(1726)));
    outputs(5432) <= (layer2_outputs(2585)) xor (layer2_outputs(2174));
    outputs(5433) <= not(layer2_outputs(158));
    outputs(5434) <= not(layer2_outputs(5992));
    outputs(5435) <= layer2_outputs(6350);
    outputs(5436) <= layer2_outputs(5115);
    outputs(5437) <= (layer2_outputs(8923)) and (layer2_outputs(6765));
    outputs(5438) <= (layer2_outputs(6184)) and (layer2_outputs(5973));
    outputs(5439) <= layer2_outputs(6986);
    outputs(5440) <= layer2_outputs(3948);
    outputs(5441) <= not(layer2_outputs(2583));
    outputs(5442) <= not(layer2_outputs(3890));
    outputs(5443) <= not(layer2_outputs(7649));
    outputs(5444) <= (layer2_outputs(3210)) and not (layer2_outputs(7066));
    outputs(5445) <= not(layer2_outputs(3583));
    outputs(5446) <= (layer2_outputs(4059)) and not (layer2_outputs(1989));
    outputs(5447) <= not(layer2_outputs(9092));
    outputs(5448) <= not((layer2_outputs(7894)) xor (layer2_outputs(2477)));
    outputs(5449) <= (layer2_outputs(9745)) xor (layer2_outputs(5296));
    outputs(5450) <= not(layer2_outputs(2350));
    outputs(5451) <= not((layer2_outputs(1615)) xor (layer2_outputs(2825)));
    outputs(5452) <= not(layer2_outputs(2727));
    outputs(5453) <= (layer2_outputs(7349)) and (layer2_outputs(1669));
    outputs(5454) <= not(layer2_outputs(3577));
    outputs(5455) <= (layer2_outputs(327)) xor (layer2_outputs(3912));
    outputs(5456) <= not(layer2_outputs(4940));
    outputs(5457) <= layer2_outputs(2381);
    outputs(5458) <= layer2_outputs(4079);
    outputs(5459) <= (layer2_outputs(2925)) and not (layer2_outputs(9794));
    outputs(5460) <= not(layer2_outputs(6219));
    outputs(5461) <= (layer2_outputs(3214)) xor (layer2_outputs(114));
    outputs(5462) <= not(layer2_outputs(8479));
    outputs(5463) <= (layer2_outputs(8034)) xor (layer2_outputs(5026));
    outputs(5464) <= not((layer2_outputs(2932)) xor (layer2_outputs(6605)));
    outputs(5465) <= not((layer2_outputs(4717)) and (layer2_outputs(2128)));
    outputs(5466) <= layer2_outputs(4678);
    outputs(5467) <= not(layer2_outputs(3253));
    outputs(5468) <= (layer2_outputs(5981)) or (layer2_outputs(1505));
    outputs(5469) <= (layer2_outputs(2750)) xor (layer2_outputs(3214));
    outputs(5470) <= layer2_outputs(5818);
    outputs(5471) <= layer2_outputs(5543);
    outputs(5472) <= (layer2_outputs(9154)) xor (layer2_outputs(6325));
    outputs(5473) <= (layer2_outputs(6666)) xor (layer2_outputs(8587));
    outputs(5474) <= layer2_outputs(8050);
    outputs(5475) <= layer2_outputs(1968);
    outputs(5476) <= layer2_outputs(8877);
    outputs(5477) <= layer2_outputs(7838);
    outputs(5478) <= not((layer2_outputs(1855)) xor (layer2_outputs(6494)));
    outputs(5479) <= (layer2_outputs(3156)) xor (layer2_outputs(6336));
    outputs(5480) <= layer2_outputs(3285);
    outputs(5481) <= not(layer2_outputs(926));
    outputs(5482) <= (layer2_outputs(4986)) and not (layer2_outputs(6073));
    outputs(5483) <= layer2_outputs(9230);
    outputs(5484) <= layer2_outputs(6022);
    outputs(5485) <= not((layer2_outputs(8136)) xor (layer2_outputs(5278)));
    outputs(5486) <= not(layer2_outputs(2483));
    outputs(5487) <= not((layer2_outputs(9276)) xor (layer2_outputs(200)));
    outputs(5488) <= (layer2_outputs(632)) and (layer2_outputs(2230));
    outputs(5489) <= not((layer2_outputs(1023)) and (layer2_outputs(2120)));
    outputs(5490) <= not(layer2_outputs(3429));
    outputs(5491) <= not(layer2_outputs(9329));
    outputs(5492) <= not((layer2_outputs(1862)) xor (layer2_outputs(3254)));
    outputs(5493) <= not(layer2_outputs(7741)) or (layer2_outputs(804));
    outputs(5494) <= layer2_outputs(5567);
    outputs(5495) <= not(layer2_outputs(3803));
    outputs(5496) <= not(layer2_outputs(4324));
    outputs(5497) <= (layer2_outputs(1560)) xor (layer2_outputs(481));
    outputs(5498) <= not(layer2_outputs(7981));
    outputs(5499) <= (layer2_outputs(3316)) and not (layer2_outputs(8448));
    outputs(5500) <= (layer2_outputs(5762)) xor (layer2_outputs(2440));
    outputs(5501) <= (layer2_outputs(9609)) xor (layer2_outputs(3859));
    outputs(5502) <= layer2_outputs(7156);
    outputs(5503) <= not(layer2_outputs(9312));
    outputs(5504) <= not(layer2_outputs(820));
    outputs(5505) <= (layer2_outputs(6816)) and not (layer2_outputs(8258));
    outputs(5506) <= not(layer2_outputs(7507)) or (layer2_outputs(9284));
    outputs(5507) <= (layer2_outputs(7495)) and not (layer2_outputs(5390));
    outputs(5508) <= not(layer2_outputs(9952));
    outputs(5509) <= not((layer2_outputs(1746)) xor (layer2_outputs(7554)));
    outputs(5510) <= layer2_outputs(8578);
    outputs(5511) <= (layer2_outputs(1224)) xor (layer2_outputs(155));
    outputs(5512) <= (layer2_outputs(853)) and (layer2_outputs(918));
    outputs(5513) <= (layer2_outputs(4427)) xor (layer2_outputs(3647));
    outputs(5514) <= not(layer2_outputs(6189));
    outputs(5515) <= (layer2_outputs(1518)) and (layer2_outputs(1448));
    outputs(5516) <= not(layer2_outputs(7543)) or (layer2_outputs(8334));
    outputs(5517) <= (layer2_outputs(7782)) xor (layer2_outputs(5179));
    outputs(5518) <= not((layer2_outputs(7328)) xor (layer2_outputs(4872)));
    outputs(5519) <= layer2_outputs(4792);
    outputs(5520) <= (layer2_outputs(1779)) and (layer2_outputs(7945));
    outputs(5521) <= (layer2_outputs(3699)) xor (layer2_outputs(48));
    outputs(5522) <= not((layer2_outputs(7178)) xor (layer2_outputs(5345)));
    outputs(5523) <= not(layer2_outputs(2380));
    outputs(5524) <= (layer2_outputs(7887)) and not (layer2_outputs(6213));
    outputs(5525) <= not((layer2_outputs(1929)) xor (layer2_outputs(6066)));
    outputs(5526) <= layer2_outputs(5602);
    outputs(5527) <= (layer2_outputs(659)) or (layer2_outputs(4133));
    outputs(5528) <= (layer2_outputs(9803)) xor (layer2_outputs(8921));
    outputs(5529) <= not(layer2_outputs(9474));
    outputs(5530) <= (layer2_outputs(1756)) xor (layer2_outputs(9237));
    outputs(5531) <= not(layer2_outputs(8806));
    outputs(5532) <= not(layer2_outputs(939));
    outputs(5533) <= not((layer2_outputs(8142)) xor (layer2_outputs(4064)));
    outputs(5534) <= layer2_outputs(4501);
    outputs(5535) <= not((layer2_outputs(2611)) or (layer2_outputs(8287)));
    outputs(5536) <= not(layer2_outputs(765));
    outputs(5537) <= not((layer2_outputs(2442)) xor (layer2_outputs(4508)));
    outputs(5538) <= not(layer2_outputs(10199));
    outputs(5539) <= not(layer2_outputs(4404));
    outputs(5540) <= layer2_outputs(9473);
    outputs(5541) <= not(layer2_outputs(106));
    outputs(5542) <= not(layer2_outputs(5172)) or (layer2_outputs(8387));
    outputs(5543) <= (layer2_outputs(3821)) xor (layer2_outputs(2150));
    outputs(5544) <= (layer2_outputs(513)) xor (layer2_outputs(1315));
    outputs(5545) <= (layer2_outputs(2344)) xor (layer2_outputs(5727));
    outputs(5546) <= not((layer2_outputs(5758)) xor (layer2_outputs(3139)));
    outputs(5547) <= layer2_outputs(883);
    outputs(5548) <= not((layer2_outputs(4244)) xor (layer2_outputs(5196)));
    outputs(5549) <= not((layer2_outputs(377)) or (layer2_outputs(8370)));
    outputs(5550) <= not(layer2_outputs(375));
    outputs(5551) <= not((layer2_outputs(2192)) and (layer2_outputs(9744)));
    outputs(5552) <= not((layer2_outputs(8464)) xor (layer2_outputs(2465)));
    outputs(5553) <= (layer2_outputs(1260)) xor (layer2_outputs(3977));
    outputs(5554) <= layer2_outputs(6303);
    outputs(5555) <= (layer2_outputs(9091)) and not (layer2_outputs(4773));
    outputs(5556) <= (layer2_outputs(2465)) xor (layer2_outputs(6152));
    outputs(5557) <= not(layer2_outputs(9773));
    outputs(5558) <= (layer2_outputs(416)) xor (layer2_outputs(9132));
    outputs(5559) <= layer2_outputs(3672);
    outputs(5560) <= not(layer2_outputs(1435)) or (layer2_outputs(6340));
    outputs(5561) <= not(layer2_outputs(2025));
    outputs(5562) <= layer2_outputs(9228);
    outputs(5563) <= not(layer2_outputs(865));
    outputs(5564) <= layer2_outputs(1684);
    outputs(5565) <= not((layer2_outputs(9093)) xor (layer2_outputs(3838)));
    outputs(5566) <= (layer2_outputs(3036)) xor (layer2_outputs(4326));
    outputs(5567) <= layer2_outputs(2688);
    outputs(5568) <= (layer2_outputs(5865)) xor (layer2_outputs(9555));
    outputs(5569) <= (layer2_outputs(8779)) xor (layer2_outputs(8896));
    outputs(5570) <= not((layer2_outputs(745)) xor (layer2_outputs(2436)));
    outputs(5571) <= not((layer2_outputs(8062)) and (layer2_outputs(3388)));
    outputs(5572) <= (layer2_outputs(3489)) xor (layer2_outputs(9095));
    outputs(5573) <= (layer2_outputs(5095)) xor (layer2_outputs(7960));
    outputs(5574) <= not((layer2_outputs(1573)) xor (layer2_outputs(1981)));
    outputs(5575) <= not(layer2_outputs(6227));
    outputs(5576) <= layer2_outputs(245);
    outputs(5577) <= not(layer2_outputs(10128));
    outputs(5578) <= not(layer2_outputs(2422));
    outputs(5579) <= not(layer2_outputs(587)) or (layer2_outputs(5618));
    outputs(5580) <= not((layer2_outputs(3939)) xor (layer2_outputs(3447)));
    outputs(5581) <= not((layer2_outputs(7612)) xor (layer2_outputs(9254)));
    outputs(5582) <= not(layer2_outputs(4591)) or (layer2_outputs(4733));
    outputs(5583) <= not(layer2_outputs(5615));
    outputs(5584) <= layer2_outputs(7723);
    outputs(5585) <= layer2_outputs(9315);
    outputs(5586) <= not((layer2_outputs(138)) xor (layer2_outputs(8102)));
    outputs(5587) <= not(layer2_outputs(198));
    outputs(5588) <= layer2_outputs(1872);
    outputs(5589) <= layer2_outputs(3132);
    outputs(5590) <= layer2_outputs(3453);
    outputs(5591) <= layer2_outputs(5154);
    outputs(5592) <= not(layer2_outputs(4639));
    outputs(5593) <= layer2_outputs(9065);
    outputs(5594) <= not(layer2_outputs(4930)) or (layer2_outputs(584));
    outputs(5595) <= not(layer2_outputs(8407));
    outputs(5596) <= layer2_outputs(1881);
    outputs(5597) <= (layer2_outputs(8299)) xor (layer2_outputs(1698));
    outputs(5598) <= layer2_outputs(2175);
    outputs(5599) <= (layer2_outputs(4355)) and (layer2_outputs(8875));
    outputs(5600) <= (layer2_outputs(154)) xor (layer2_outputs(2747));
    outputs(5601) <= layer2_outputs(5570);
    outputs(5602) <= layer2_outputs(8233);
    outputs(5603) <= layer2_outputs(934);
    outputs(5604) <= layer2_outputs(9205);
    outputs(5605) <= not(layer2_outputs(6024));
    outputs(5606) <= not(layer2_outputs(2775));
    outputs(5607) <= not(layer2_outputs(10191));
    outputs(5608) <= layer2_outputs(8477);
    outputs(5609) <= (layer2_outputs(6385)) xor (layer2_outputs(9680));
    outputs(5610) <= not(layer2_outputs(2245));
    outputs(5611) <= not((layer2_outputs(3773)) xor (layer2_outputs(7228)));
    outputs(5612) <= not((layer2_outputs(1101)) xor (layer2_outputs(2781)));
    outputs(5613) <= layer2_outputs(6306);
    outputs(5614) <= (layer2_outputs(7275)) and (layer2_outputs(460));
    outputs(5615) <= (layer2_outputs(6125)) xor (layer2_outputs(6021));
    outputs(5616) <= (layer2_outputs(4126)) and not (layer2_outputs(5624));
    outputs(5617) <= layer2_outputs(6446);
    outputs(5618) <= layer2_outputs(2929);
    outputs(5619) <= (layer2_outputs(9657)) xor (layer2_outputs(695));
    outputs(5620) <= not((layer2_outputs(5451)) xor (layer2_outputs(2088)));
    outputs(5621) <= not(layer2_outputs(7714));
    outputs(5622) <= (layer2_outputs(2254)) and not (layer2_outputs(1806));
    outputs(5623) <= not(layer2_outputs(1216));
    outputs(5624) <= layer2_outputs(2629);
    outputs(5625) <= layer2_outputs(7182);
    outputs(5626) <= (layer2_outputs(7114)) xor (layer2_outputs(6666));
    outputs(5627) <= not(layer2_outputs(1308));
    outputs(5628) <= not((layer2_outputs(8480)) xor (layer2_outputs(6726)));
    outputs(5629) <= not((layer2_outputs(4748)) or (layer2_outputs(4006)));
    outputs(5630) <= layer2_outputs(4197);
    outputs(5631) <= layer2_outputs(3353);
    outputs(5632) <= not(layer2_outputs(3498));
    outputs(5633) <= (layer2_outputs(4848)) xor (layer2_outputs(7523));
    outputs(5634) <= not((layer2_outputs(9256)) xor (layer2_outputs(9980)));
    outputs(5635) <= layer2_outputs(7574);
    outputs(5636) <= not(layer2_outputs(4166)) or (layer2_outputs(4361));
    outputs(5637) <= not(layer2_outputs(2489)) or (layer2_outputs(8904));
    outputs(5638) <= not((layer2_outputs(1317)) xor (layer2_outputs(8301)));
    outputs(5639) <= not(layer2_outputs(7318));
    outputs(5640) <= not(layer2_outputs(3611));
    outputs(5641) <= layer2_outputs(3809);
    outputs(5642) <= not((layer2_outputs(8989)) or (layer2_outputs(583)));
    outputs(5643) <= not((layer2_outputs(4182)) xor (layer2_outputs(3384)));
    outputs(5644) <= layer2_outputs(567);
    outputs(5645) <= layer2_outputs(4644);
    outputs(5646) <= not(layer2_outputs(4303));
    outputs(5647) <= not(layer2_outputs(7984));
    outputs(5648) <= not((layer2_outputs(6086)) and (layer2_outputs(6324)));
    outputs(5649) <= layer2_outputs(5054);
    outputs(5650) <= (layer2_outputs(2884)) and (layer2_outputs(9880));
    outputs(5651) <= layer2_outputs(2692);
    outputs(5652) <= (layer2_outputs(2927)) xor (layer2_outputs(36));
    outputs(5653) <= layer2_outputs(9377);
    outputs(5654) <= layer2_outputs(7911);
    outputs(5655) <= not((layer2_outputs(5815)) and (layer2_outputs(1019)));
    outputs(5656) <= layer2_outputs(3663);
    outputs(5657) <= not(layer2_outputs(8993));
    outputs(5658) <= not(layer2_outputs(7137));
    outputs(5659) <= layer2_outputs(846);
    outputs(5660) <= not((layer2_outputs(9038)) or (layer2_outputs(3749)));
    outputs(5661) <= not((layer2_outputs(4827)) or (layer2_outputs(8725)));
    outputs(5662) <= layer2_outputs(4079);
    outputs(5663) <= (layer2_outputs(21)) and not (layer2_outputs(9558));
    outputs(5664) <= layer2_outputs(4742);
    outputs(5665) <= layer2_outputs(3779);
    outputs(5666) <= (layer2_outputs(1614)) xor (layer2_outputs(4526));
    outputs(5667) <= not(layer2_outputs(2151));
    outputs(5668) <= (layer2_outputs(3814)) xor (layer2_outputs(6483));
    outputs(5669) <= (layer2_outputs(2079)) xor (layer2_outputs(237));
    outputs(5670) <= not((layer2_outputs(8822)) xor (layer2_outputs(4480)));
    outputs(5671) <= not(layer2_outputs(2103)) or (layer2_outputs(892));
    outputs(5672) <= not((layer2_outputs(3950)) xor (layer2_outputs(4484)));
    outputs(5673) <= not((layer2_outputs(76)) xor (layer2_outputs(6767)));
    outputs(5674) <= layer2_outputs(3641);
    outputs(5675) <= (layer2_outputs(5056)) xor (layer2_outputs(8432));
    outputs(5676) <= (layer2_outputs(698)) xor (layer2_outputs(416));
    outputs(5677) <= not(layer2_outputs(2244));
    outputs(5678) <= not((layer2_outputs(5105)) or (layer2_outputs(5373)));
    outputs(5679) <= layer2_outputs(6022);
    outputs(5680) <= layer2_outputs(6939);
    outputs(5681) <= (layer2_outputs(3760)) xor (layer2_outputs(1381));
    outputs(5682) <= not(layer2_outputs(226));
    outputs(5683) <= (layer2_outputs(6419)) xor (layer2_outputs(2326));
    outputs(5684) <= not((layer2_outputs(1780)) or (layer2_outputs(9768)));
    outputs(5685) <= not((layer2_outputs(7237)) xor (layer2_outputs(203)));
    outputs(5686) <= (layer2_outputs(5990)) and not (layer2_outputs(2907));
    outputs(5687) <= not(layer2_outputs(6238)) or (layer2_outputs(589));
    outputs(5688) <= not(layer2_outputs(8593));
    outputs(5689) <= layer2_outputs(6093);
    outputs(5690) <= layer2_outputs(2399);
    outputs(5691) <= not(layer2_outputs(7273));
    outputs(5692) <= not((layer2_outputs(6358)) xor (layer2_outputs(7560)));
    outputs(5693) <= not(layer2_outputs(9700)) or (layer2_outputs(3900));
    outputs(5694) <= not(layer2_outputs(4156));
    outputs(5695) <= not((layer2_outputs(8461)) xor (layer2_outputs(5437)));
    outputs(5696) <= layer2_outputs(2078);
    outputs(5697) <= layer2_outputs(1586);
    outputs(5698) <= (layer2_outputs(5882)) xor (layer2_outputs(1195));
    outputs(5699) <= not(layer2_outputs(1013)) or (layer2_outputs(9397));
    outputs(5700) <= not(layer2_outputs(6570));
    outputs(5701) <= not(layer2_outputs(7951));
    outputs(5702) <= not(layer2_outputs(1166));
    outputs(5703) <= not(layer2_outputs(4404));
    outputs(5704) <= layer2_outputs(9895);
    outputs(5705) <= (layer2_outputs(1442)) xor (layer2_outputs(1930));
    outputs(5706) <= not(layer2_outputs(8350));
    outputs(5707) <= not((layer2_outputs(8326)) xor (layer2_outputs(7722)));
    outputs(5708) <= (layer2_outputs(7772)) and not (layer2_outputs(9296));
    outputs(5709) <= not(layer2_outputs(2210));
    outputs(5710) <= layer2_outputs(9335);
    outputs(5711) <= not(layer2_outputs(1318));
    outputs(5712) <= layer2_outputs(212);
    outputs(5713) <= layer2_outputs(1775);
    outputs(5714) <= layer2_outputs(2876);
    outputs(5715) <= layer2_outputs(2681);
    outputs(5716) <= (layer2_outputs(5153)) and not (layer2_outputs(2160));
    outputs(5717) <= (layer2_outputs(5847)) and not (layer2_outputs(9499));
    outputs(5718) <= not(layer2_outputs(1629));
    outputs(5719) <= not((layer2_outputs(1862)) xor (layer2_outputs(7676)));
    outputs(5720) <= (layer2_outputs(7846)) xor (layer2_outputs(1418));
    outputs(5721) <= not((layer2_outputs(7179)) xor (layer2_outputs(3092)));
    outputs(5722) <= not((layer2_outputs(805)) xor (layer2_outputs(9350)));
    outputs(5723) <= (layer2_outputs(2515)) and not (layer2_outputs(2780));
    outputs(5724) <= not(layer2_outputs(7557));
    outputs(5725) <= not((layer2_outputs(5596)) xor (layer2_outputs(2817)));
    outputs(5726) <= not(layer2_outputs(9836));
    outputs(5727) <= not(layer2_outputs(2731));
    outputs(5728) <= (layer2_outputs(6252)) xor (layer2_outputs(10089));
    outputs(5729) <= layer2_outputs(3315);
    outputs(5730) <= layer2_outputs(3244);
    outputs(5731) <= layer2_outputs(6801);
    outputs(5732) <= layer2_outputs(6544);
    outputs(5733) <= not(layer2_outputs(5244)) or (layer2_outputs(1875));
    outputs(5734) <= not(layer2_outputs(1976));
    outputs(5735) <= layer2_outputs(821);
    outputs(5736) <= not((layer2_outputs(3418)) xor (layer2_outputs(891)));
    outputs(5737) <= layer2_outputs(8249);
    outputs(5738) <= (layer2_outputs(1066)) xor (layer2_outputs(7759));
    outputs(5739) <= not((layer2_outputs(8141)) xor (layer2_outputs(2607)));
    outputs(5740) <= (layer2_outputs(9658)) and (layer2_outputs(3716));
    outputs(5741) <= layer2_outputs(834);
    outputs(5742) <= not(layer2_outputs(3166));
    outputs(5743) <= not(layer2_outputs(4542));
    outputs(5744) <= not(layer2_outputs(3786));
    outputs(5745) <= (layer2_outputs(7758)) xor (layer2_outputs(5827));
    outputs(5746) <= not(layer2_outputs(3903));
    outputs(5747) <= not(layer2_outputs(1576)) or (layer2_outputs(7881));
    outputs(5748) <= (layer2_outputs(9761)) and not (layer2_outputs(3001));
    outputs(5749) <= layer2_outputs(5386);
    outputs(5750) <= not(layer2_outputs(10056));
    outputs(5751) <= layer2_outputs(5610);
    outputs(5752) <= layer2_outputs(5796);
    outputs(5753) <= layer2_outputs(5595);
    outputs(5754) <= (layer2_outputs(928)) xor (layer2_outputs(5848));
    outputs(5755) <= not(layer2_outputs(3881));
    outputs(5756) <= layer2_outputs(5221);
    outputs(5757) <= layer2_outputs(2955);
    outputs(5758) <= layer2_outputs(8321);
    outputs(5759) <= not(layer2_outputs(4496));
    outputs(5760) <= (layer2_outputs(8474)) xor (layer2_outputs(1159));
    outputs(5761) <= (layer2_outputs(8439)) xor (layer2_outputs(9225));
    outputs(5762) <= not((layer2_outputs(1514)) or (layer2_outputs(1932)));
    outputs(5763) <= not((layer2_outputs(9951)) and (layer2_outputs(6046)));
    outputs(5764) <= (layer2_outputs(3679)) xor (layer2_outputs(7617));
    outputs(5765) <= layer2_outputs(3060);
    outputs(5766) <= layer2_outputs(3107);
    outputs(5767) <= layer2_outputs(4229);
    outputs(5768) <= (layer2_outputs(7053)) xor (layer2_outputs(3805));
    outputs(5769) <= layer2_outputs(9426);
    outputs(5770) <= not(layer2_outputs(2307)) or (layer2_outputs(731));
    outputs(5771) <= (layer2_outputs(6154)) xor (layer2_outputs(5382));
    outputs(5772) <= not(layer2_outputs(5633));
    outputs(5773) <= (layer2_outputs(8678)) xor (layer2_outputs(5654));
    outputs(5774) <= (layer2_outputs(9083)) xor (layer2_outputs(8430));
    outputs(5775) <= not(layer2_outputs(2872));
    outputs(5776) <= (layer2_outputs(5250)) xor (layer2_outputs(4106));
    outputs(5777) <= (layer2_outputs(9253)) xor (layer2_outputs(699));
    outputs(5778) <= layer2_outputs(851);
    outputs(5779) <= layer2_outputs(2634);
    outputs(5780) <= not(layer2_outputs(6063));
    outputs(5781) <= not(layer2_outputs(3796)) or (layer2_outputs(1332));
    outputs(5782) <= not(layer2_outputs(4524));
    outputs(5783) <= not(layer2_outputs(4567));
    outputs(5784) <= (layer2_outputs(295)) xor (layer2_outputs(1894));
    outputs(5785) <= layer2_outputs(8068);
    outputs(5786) <= (layer2_outputs(660)) xor (layer2_outputs(5280));
    outputs(5787) <= not((layer2_outputs(10143)) or (layer2_outputs(4663)));
    outputs(5788) <= (layer2_outputs(6533)) or (layer2_outputs(4665));
    outputs(5789) <= not((layer2_outputs(8446)) xor (layer2_outputs(5184)));
    outputs(5790) <= not(layer2_outputs(3461));
    outputs(5791) <= not((layer2_outputs(6445)) xor (layer2_outputs(6303)));
    outputs(5792) <= layer2_outputs(8659);
    outputs(5793) <= not(layer2_outputs(6923));
    outputs(5794) <= (layer2_outputs(6175)) and not (layer2_outputs(4516));
    outputs(5795) <= not(layer2_outputs(6311));
    outputs(5796) <= not(layer2_outputs(5226));
    outputs(5797) <= (layer2_outputs(7038)) and not (layer2_outputs(9853));
    outputs(5798) <= not((layer2_outputs(1940)) xor (layer2_outputs(2793)));
    outputs(5799) <= (layer2_outputs(9308)) xor (layer2_outputs(8045));
    outputs(5800) <= (layer2_outputs(4024)) xor (layer2_outputs(9716));
    outputs(5801) <= (layer2_outputs(2267)) and not (layer2_outputs(3688));
    outputs(5802) <= not(layer2_outputs(1027));
    outputs(5803) <= (layer2_outputs(3121)) xor (layer2_outputs(6463));
    outputs(5804) <= not(layer2_outputs(8168));
    outputs(5805) <= not(layer2_outputs(1478)) or (layer2_outputs(9457));
    outputs(5806) <= not(layer2_outputs(8270));
    outputs(5807) <= (layer2_outputs(4116)) and (layer2_outputs(9567));
    outputs(5808) <= not(layer2_outputs(3838));
    outputs(5809) <= (layer2_outputs(682)) and not (layer2_outputs(664));
    outputs(5810) <= layer2_outputs(2698);
    outputs(5811) <= not(layer2_outputs(6300));
    outputs(5812) <= (layer2_outputs(6852)) and (layer2_outputs(3473));
    outputs(5813) <= not(layer2_outputs(765));
    outputs(5814) <= layer2_outputs(2698);
    outputs(5815) <= not(layer2_outputs(163)) or (layer2_outputs(3888));
    outputs(5816) <= not((layer2_outputs(4942)) xor (layer2_outputs(5573)));
    outputs(5817) <= not((layer2_outputs(9891)) xor (layer2_outputs(2102)));
    outputs(5818) <= layer2_outputs(7561);
    outputs(5819) <= layer2_outputs(392);
    outputs(5820) <= not((layer2_outputs(523)) xor (layer2_outputs(4611)));
    outputs(5821) <= not(layer2_outputs(6227));
    outputs(5822) <= (layer2_outputs(3072)) and not (layer2_outputs(5819));
    outputs(5823) <= not(layer2_outputs(2438));
    outputs(5824) <= not(layer2_outputs(7272));
    outputs(5825) <= layer2_outputs(6781);
    outputs(5826) <= not(layer2_outputs(907));
    outputs(5827) <= not((layer2_outputs(1722)) xor (layer2_outputs(7922)));
    outputs(5828) <= layer2_outputs(2357);
    outputs(5829) <= not((layer2_outputs(1790)) xor (layer2_outputs(8729)));
    outputs(5830) <= layer2_outputs(4193);
    outputs(5831) <= layer2_outputs(8961);
    outputs(5832) <= layer2_outputs(149);
    outputs(5833) <= not((layer2_outputs(2965)) and (layer2_outputs(5861)));
    outputs(5834) <= (layer2_outputs(5886)) xor (layer2_outputs(5856));
    outputs(5835) <= not((layer2_outputs(850)) or (layer2_outputs(5021)));
    outputs(5836) <= (layer2_outputs(1371)) and not (layer2_outputs(6198));
    outputs(5837) <= (layer2_outputs(6258)) and not (layer2_outputs(8534));
    outputs(5838) <= (layer2_outputs(5682)) and (layer2_outputs(3905));
    outputs(5839) <= layer2_outputs(9683);
    outputs(5840) <= (layer2_outputs(1724)) and not (layer2_outputs(2498));
    outputs(5841) <= not(layer2_outputs(5687)) or (layer2_outputs(5842));
    outputs(5842) <= not((layer2_outputs(7393)) and (layer2_outputs(5962)));
    outputs(5843) <= layer2_outputs(2535);
    outputs(5844) <= not(layer2_outputs(5082));
    outputs(5845) <= layer2_outputs(4213);
    outputs(5846) <= layer2_outputs(3979);
    outputs(5847) <= layer2_outputs(7440);
    outputs(5848) <= layer2_outputs(4753);
    outputs(5849) <= not(layer2_outputs(3064));
    outputs(5850) <= layer2_outputs(7772);
    outputs(5851) <= (layer2_outputs(8304)) and not (layer2_outputs(6856));
    outputs(5852) <= (layer2_outputs(31)) xor (layer2_outputs(5790));
    outputs(5853) <= layer2_outputs(9955);
    outputs(5854) <= layer2_outputs(8779);
    outputs(5855) <= (layer2_outputs(6494)) xor (layer2_outputs(5966));
    outputs(5856) <= layer2_outputs(2703);
    outputs(5857) <= layer2_outputs(5764);
    outputs(5858) <= not(layer2_outputs(8674));
    outputs(5859) <= layer2_outputs(9978);
    outputs(5860) <= layer2_outputs(4020);
    outputs(5861) <= (layer2_outputs(4499)) or (layer2_outputs(6761));
    outputs(5862) <= not(layer2_outputs(8038));
    outputs(5863) <= (layer2_outputs(1823)) xor (layer2_outputs(4875));
    outputs(5864) <= layer2_outputs(8320);
    outputs(5865) <= (layer2_outputs(9715)) xor (layer2_outputs(8510));
    outputs(5866) <= not(layer2_outputs(4881));
    outputs(5867) <= layer2_outputs(6061);
    outputs(5868) <= not(layer2_outputs(4776));
    outputs(5869) <= layer2_outputs(1394);
    outputs(5870) <= (layer2_outputs(7376)) xor (layer2_outputs(1356));
    outputs(5871) <= not((layer2_outputs(7366)) xor (layer2_outputs(10220)));
    outputs(5872) <= not((layer2_outputs(8178)) and (layer2_outputs(2365)));
    outputs(5873) <= layer2_outputs(8985);
    outputs(5874) <= not((layer2_outputs(9058)) xor (layer2_outputs(2232)));
    outputs(5875) <= (layer2_outputs(3471)) and (layer2_outputs(1104));
    outputs(5876) <= not((layer2_outputs(7638)) xor (layer2_outputs(4281)));
    outputs(5877) <= not((layer2_outputs(5475)) or (layer2_outputs(2305)));
    outputs(5878) <= (layer2_outputs(5991)) xor (layer2_outputs(8628));
    outputs(5879) <= not((layer2_outputs(1314)) xor (layer2_outputs(1221)));
    outputs(5880) <= not((layer2_outputs(7899)) xor (layer2_outputs(2149)));
    outputs(5881) <= not((layer2_outputs(4050)) xor (layer2_outputs(1740)));
    outputs(5882) <= not(layer2_outputs(8285));
    outputs(5883) <= layer2_outputs(1453);
    outputs(5884) <= layer2_outputs(3543);
    outputs(5885) <= not((layer2_outputs(4699)) xor (layer2_outputs(673)));
    outputs(5886) <= layer2_outputs(2369);
    outputs(5887) <= not(layer2_outputs(5992));
    outputs(5888) <= layer2_outputs(653);
    outputs(5889) <= not(layer2_outputs(8226));
    outputs(5890) <= layer2_outputs(10228);
    outputs(5891) <= not(layer2_outputs(10040));
    outputs(5892) <= not(layer2_outputs(8154));
    outputs(5893) <= not((layer2_outputs(2947)) xor (layer2_outputs(767)));
    outputs(5894) <= (layer2_outputs(4723)) xor (layer2_outputs(2946));
    outputs(5895) <= not(layer2_outputs(9773));
    outputs(5896) <= not(layer2_outputs(2527));
    outputs(5897) <= not(layer2_outputs(9463));
    outputs(5898) <= layer2_outputs(4745);
    outputs(5899) <= not(layer2_outputs(3091));
    outputs(5900) <= layer2_outputs(5572);
    outputs(5901) <= not(layer2_outputs(6788));
    outputs(5902) <= not((layer2_outputs(9277)) and (layer2_outputs(1611)));
    outputs(5903) <= layer2_outputs(8588);
    outputs(5904) <= (layer2_outputs(8518)) or (layer2_outputs(3586));
    outputs(5905) <= layer2_outputs(3033);
    outputs(5906) <= not((layer2_outputs(71)) xor (layer2_outputs(415)));
    outputs(5907) <= not(layer2_outputs(3759));
    outputs(5908) <= (layer2_outputs(7259)) xor (layer2_outputs(6055));
    outputs(5909) <= (layer2_outputs(2836)) xor (layer2_outputs(4097));
    outputs(5910) <= not((layer2_outputs(553)) xor (layer2_outputs(2379)));
    outputs(5911) <= not(layer2_outputs(8350));
    outputs(5912) <= (layer2_outputs(8746)) xor (layer2_outputs(1522));
    outputs(5913) <= layer2_outputs(7302);
    outputs(5914) <= not((layer2_outputs(6728)) or (layer2_outputs(8409)));
    outputs(5915) <= layer2_outputs(8817);
    outputs(5916) <= (layer2_outputs(3642)) xor (layer2_outputs(5504));
    outputs(5917) <= not((layer2_outputs(9832)) xor (layer2_outputs(9776)));
    outputs(5918) <= (layer2_outputs(7104)) xor (layer2_outputs(98));
    outputs(5919) <= not((layer2_outputs(1652)) xor (layer2_outputs(8783)));
    outputs(5920) <= not(layer2_outputs(304));
    outputs(5921) <= not((layer2_outputs(9738)) or (layer2_outputs(3459)));
    outputs(5922) <= not(layer2_outputs(781));
    outputs(5923) <= layer2_outputs(2230);
    outputs(5924) <= not(layer2_outputs(4232));
    outputs(5925) <= (layer2_outputs(9969)) and not (layer2_outputs(2124));
    outputs(5926) <= not(layer2_outputs(6305));
    outputs(5927) <= not(layer2_outputs(2567)) or (layer2_outputs(5272));
    outputs(5928) <= not((layer2_outputs(3670)) xor (layer2_outputs(6529)));
    outputs(5929) <= not((layer2_outputs(249)) xor (layer2_outputs(9241)));
    outputs(5930) <= not(layer2_outputs(1452));
    outputs(5931) <= not(layer2_outputs(2349));
    outputs(5932) <= not(layer2_outputs(1390));
    outputs(5933) <= not((layer2_outputs(4334)) xor (layer2_outputs(1254)));
    outputs(5934) <= layer2_outputs(6017);
    outputs(5935) <= layer2_outputs(7656);
    outputs(5936) <= layer2_outputs(6413);
    outputs(5937) <= not(layer2_outputs(8990));
    outputs(5938) <= (layer2_outputs(2997)) xor (layer2_outputs(7197));
    outputs(5939) <= not(layer2_outputs(2877));
    outputs(5940) <= (layer2_outputs(8040)) and not (layer2_outputs(5683));
    outputs(5941) <= not(layer2_outputs(7908)) or (layer2_outputs(1351));
    outputs(5942) <= layer2_outputs(2954);
    outputs(5943) <= not(layer2_outputs(6653));
    outputs(5944) <= (layer2_outputs(4788)) xor (layer2_outputs(3934));
    outputs(5945) <= layer2_outputs(1589);
    outputs(5946) <= (layer2_outputs(7763)) xor (layer2_outputs(2654));
    outputs(5947) <= layer2_outputs(4505);
    outputs(5948) <= (layer2_outputs(6280)) xor (layer2_outputs(9114));
    outputs(5949) <= layer2_outputs(9278);
    outputs(5950) <= layer2_outputs(9521);
    outputs(5951) <= not(layer2_outputs(8287));
    outputs(5952) <= not(layer2_outputs(9086));
    outputs(5953) <= not(layer2_outputs(4290)) or (layer2_outputs(9694));
    outputs(5954) <= layer2_outputs(1292);
    outputs(5955) <= layer2_outputs(1724);
    outputs(5956) <= not((layer2_outputs(1281)) and (layer2_outputs(3901)));
    outputs(5957) <= layer2_outputs(5312);
    outputs(5958) <= not((layer2_outputs(1087)) xor (layer2_outputs(4186)));
    outputs(5959) <= (layer2_outputs(4783)) and not (layer2_outputs(3953));
    outputs(5960) <= layer2_outputs(5281);
    outputs(5961) <= not(layer2_outputs(9484));
    outputs(5962) <= not((layer2_outputs(2617)) xor (layer2_outputs(4955)));
    outputs(5963) <= not(layer2_outputs(5033));
    outputs(5964) <= layer2_outputs(860);
    outputs(5965) <= (layer2_outputs(4581)) xor (layer2_outputs(1073));
    outputs(5966) <= layer2_outputs(3655);
    outputs(5967) <= (layer2_outputs(3233)) and not (layer2_outputs(7540));
    outputs(5968) <= (layer2_outputs(9658)) xor (layer2_outputs(6669));
    outputs(5969) <= not(layer2_outputs(3726));
    outputs(5970) <= not((layer2_outputs(8944)) and (layer2_outputs(2511)));
    outputs(5971) <= not((layer2_outputs(8095)) xor (layer2_outputs(7509)));
    outputs(5972) <= (layer2_outputs(6218)) and not (layer2_outputs(2686));
    outputs(5973) <= layer2_outputs(4927);
    outputs(5974) <= not(layer2_outputs(9324));
    outputs(5975) <= layer2_outputs(6523);
    outputs(5976) <= not((layer2_outputs(8383)) and (layer2_outputs(1720)));
    outputs(5977) <= (layer2_outputs(9273)) and not (layer2_outputs(9286));
    outputs(5978) <= (layer2_outputs(4244)) xor (layer2_outputs(6005));
    outputs(5979) <= layer2_outputs(7521);
    outputs(5980) <= not((layer2_outputs(8727)) or (layer2_outputs(6689)));
    outputs(5981) <= not((layer2_outputs(8421)) and (layer2_outputs(1503)));
    outputs(5982) <= not((layer2_outputs(2835)) xor (layer2_outputs(1206)));
    outputs(5983) <= layer2_outputs(8558);
    outputs(5984) <= not((layer2_outputs(438)) xor (layer2_outputs(2875)));
    outputs(5985) <= not(layer2_outputs(7921));
    outputs(5986) <= not(layer2_outputs(1204));
    outputs(5987) <= not((layer2_outputs(5041)) xor (layer2_outputs(8925)));
    outputs(5988) <= (layer2_outputs(8684)) and not (layer2_outputs(8739));
    outputs(5989) <= layer2_outputs(10080);
    outputs(5990) <= not((layer2_outputs(7694)) xor (layer2_outputs(4337)));
    outputs(5991) <= (layer2_outputs(6743)) and not (layer2_outputs(3659));
    outputs(5992) <= not((layer2_outputs(2974)) xor (layer2_outputs(9867)));
    outputs(5993) <= (layer2_outputs(2444)) xor (layer2_outputs(4886));
    outputs(5994) <= (layer2_outputs(7120)) xor (layer2_outputs(3546));
    outputs(5995) <= not((layer2_outputs(7813)) xor (layer2_outputs(5852)));
    outputs(5996) <= layer2_outputs(6951);
    outputs(5997) <= not((layer2_outputs(4517)) xor (layer2_outputs(7360)));
    outputs(5998) <= not((layer2_outputs(6287)) xor (layer2_outputs(1088)));
    outputs(5999) <= layer2_outputs(6810);
    outputs(6000) <= (layer2_outputs(6853)) and (layer2_outputs(2910));
    outputs(6001) <= layer2_outputs(2213);
    outputs(6002) <= layer2_outputs(5296);
    outputs(6003) <= layer2_outputs(7814);
    outputs(6004) <= (layer2_outputs(7206)) and not (layer2_outputs(6556));
    outputs(6005) <= not(layer2_outputs(9164));
    outputs(6006) <= not((layer2_outputs(6120)) and (layer2_outputs(1765)));
    outputs(6007) <= layer2_outputs(3795);
    outputs(6008) <= (layer2_outputs(850)) xor (layer2_outputs(8636));
    outputs(6009) <= (layer2_outputs(3502)) and not (layer2_outputs(9113));
    outputs(6010) <= (layer2_outputs(9023)) xor (layer2_outputs(8542));
    outputs(6011) <= not(layer2_outputs(7806)) or (layer2_outputs(835));
    outputs(6012) <= not(layer2_outputs(7573));
    outputs(6013) <= not(layer2_outputs(8736));
    outputs(6014) <= not((layer2_outputs(8046)) xor (layer2_outputs(5874)));
    outputs(6015) <= layer2_outputs(3085);
    outputs(6016) <= (layer2_outputs(7336)) and (layer2_outputs(5107));
    outputs(6017) <= layer2_outputs(4072);
    outputs(6018) <= (layer2_outputs(8975)) xor (layer2_outputs(473));
    outputs(6019) <= not((layer2_outputs(9383)) xor (layer2_outputs(2513)));
    outputs(6020) <= not((layer2_outputs(2429)) xor (layer2_outputs(10152)));
    outputs(6021) <= (layer2_outputs(111)) xor (layer2_outputs(234));
    outputs(6022) <= not(layer2_outputs(7162));
    outputs(6023) <= layer2_outputs(1191);
    outputs(6024) <= not(layer2_outputs(8869));
    outputs(6025) <= not((layer2_outputs(565)) xor (layer2_outputs(1169)));
    outputs(6026) <= layer2_outputs(9567);
    outputs(6027) <= not(layer2_outputs(2447)) or (layer2_outputs(4975));
    outputs(6028) <= not(layer2_outputs(3154));
    outputs(6029) <= (layer2_outputs(3624)) and not (layer2_outputs(3665));
    outputs(6030) <= layer2_outputs(5952);
    outputs(6031) <= (layer2_outputs(2800)) xor (layer2_outputs(9829));
    outputs(6032) <= not(layer2_outputs(6260));
    outputs(6033) <= (layer2_outputs(9163)) xor (layer2_outputs(4289));
    outputs(6034) <= (layer2_outputs(3428)) and not (layer2_outputs(9681));
    outputs(6035) <= layer2_outputs(6852);
    outputs(6036) <= not(layer2_outputs(10226));
    outputs(6037) <= (layer2_outputs(6581)) and not (layer2_outputs(2144));
    outputs(6038) <= not(layer2_outputs(2227));
    outputs(6039) <= not((layer2_outputs(6378)) xor (layer2_outputs(8869)));
    outputs(6040) <= (layer2_outputs(5575)) or (layer2_outputs(3021));
    outputs(6041) <= not((layer2_outputs(789)) xor (layer2_outputs(3199)));
    outputs(6042) <= layer2_outputs(7107);
    outputs(6043) <= not((layer2_outputs(9636)) xor (layer2_outputs(2169)));
    outputs(6044) <= not(layer2_outputs(385)) or (layer2_outputs(9425));
    outputs(6045) <= layer2_outputs(8918);
    outputs(6046) <= not((layer2_outputs(4388)) xor (layer2_outputs(7550)));
    outputs(6047) <= not((layer2_outputs(961)) xor (layer2_outputs(7506)));
    outputs(6048) <= not(layer2_outputs(102));
    outputs(6049) <= layer2_outputs(3927);
    outputs(6050) <= layer2_outputs(3928);
    outputs(6051) <= not((layer2_outputs(8131)) xor (layer2_outputs(1666)));
    outputs(6052) <= layer2_outputs(4126);
    outputs(6053) <= not(layer2_outputs(2721));
    outputs(6054) <= not(layer2_outputs(5787));
    outputs(6055) <= layer2_outputs(7835);
    outputs(6056) <= not((layer2_outputs(240)) and (layer2_outputs(1671)));
    outputs(6057) <= layer2_outputs(7334);
    outputs(6058) <= layer2_outputs(9974);
    outputs(6059) <= (layer2_outputs(1627)) xor (layer2_outputs(4209));
    outputs(6060) <= not((layer2_outputs(5849)) xor (layer2_outputs(4635)));
    outputs(6061) <= (layer2_outputs(4268)) xor (layer2_outputs(7142));
    outputs(6062) <= not((layer2_outputs(4219)) xor (layer2_outputs(8016)));
    outputs(6063) <= layer2_outputs(2153);
    outputs(6064) <= (layer2_outputs(46)) and (layer2_outputs(10041));
    outputs(6065) <= layer2_outputs(1071);
    outputs(6066) <= not(layer2_outputs(5101));
    outputs(6067) <= layer2_outputs(5334);
    outputs(6068) <= not((layer2_outputs(679)) xor (layer2_outputs(4187)));
    outputs(6069) <= (layer2_outputs(189)) and (layer2_outputs(460));
    outputs(6070) <= not(layer2_outputs(9309));
    outputs(6071) <= not(layer2_outputs(1137));
    outputs(6072) <= not(layer2_outputs(594));
    outputs(6073) <= (layer2_outputs(2848)) xor (layer2_outputs(4966));
    outputs(6074) <= not((layer2_outputs(7748)) or (layer2_outputs(757)));
    outputs(6075) <= layer2_outputs(2950);
    outputs(6076) <= not((layer2_outputs(4643)) xor (layer2_outputs(9093)));
    outputs(6077) <= (layer2_outputs(8490)) xor (layer2_outputs(8176));
    outputs(6078) <= not(layer2_outputs(5801));
    outputs(6079) <= not(layer2_outputs(1942)) or (layer2_outputs(7339));
    outputs(6080) <= not((layer2_outputs(4082)) or (layer2_outputs(3043)));
    outputs(6081) <= not((layer2_outputs(4542)) and (layer2_outputs(242)));
    outputs(6082) <= (layer2_outputs(5599)) xor (layer2_outputs(7118));
    outputs(6083) <= not(layer2_outputs(8897));
    outputs(6084) <= (layer2_outputs(6429)) and not (layer2_outputs(3098));
    outputs(6085) <= not((layer2_outputs(6637)) xor (layer2_outputs(2945)));
    outputs(6086) <= not((layer2_outputs(4168)) xor (layer2_outputs(279)));
    outputs(6087) <= not(layer2_outputs(1208));
    outputs(6088) <= not((layer2_outputs(3496)) xor (layer2_outputs(2372)));
    outputs(6089) <= (layer2_outputs(9889)) xor (layer2_outputs(7452));
    outputs(6090) <= (layer2_outputs(8958)) xor (layer2_outputs(1967));
    outputs(6091) <= not(layer2_outputs(2701));
    outputs(6092) <= not((layer2_outputs(1202)) xor (layer2_outputs(3967)));
    outputs(6093) <= not(layer2_outputs(4510));
    outputs(6094) <= not((layer2_outputs(3785)) xor (layer2_outputs(8744)));
    outputs(6095) <= not(layer2_outputs(7876));
    outputs(6096) <= layer2_outputs(5034);
    outputs(6097) <= layer2_outputs(2925);
    outputs(6098) <= not(layer2_outputs(7177));
    outputs(6099) <= not((layer2_outputs(9020)) xor (layer2_outputs(73)));
    outputs(6100) <= not(layer2_outputs(2105));
    outputs(6101) <= layer2_outputs(2014);
    outputs(6102) <= layer2_outputs(8652);
    outputs(6103) <= (layer2_outputs(3330)) xor (layer2_outputs(6088));
    outputs(6104) <= (layer2_outputs(1776)) xor (layer2_outputs(1141));
    outputs(6105) <= (layer2_outputs(6872)) xor (layer2_outputs(2660));
    outputs(6106) <= not(layer2_outputs(2359));
    outputs(6107) <= not(layer2_outputs(1923));
    outputs(6108) <= not(layer2_outputs(3855));
    outputs(6109) <= not(layer2_outputs(8871));
    outputs(6110) <= layer2_outputs(6162);
    outputs(6111) <= not(layer2_outputs(4418));
    outputs(6112) <= layer2_outputs(693);
    outputs(6113) <= (layer2_outputs(10179)) xor (layer2_outputs(386));
    outputs(6114) <= not(layer2_outputs(8060));
    outputs(6115) <= layer2_outputs(7696);
    outputs(6116) <= not(layer2_outputs(9763));
    outputs(6117) <= not((layer2_outputs(4702)) xor (layer2_outputs(9285)));
    outputs(6118) <= layer2_outputs(10001);
    outputs(6119) <= not(layer2_outputs(5553)) or (layer2_outputs(9582));
    outputs(6120) <= not(layer2_outputs(3153));
    outputs(6121) <= not((layer2_outputs(677)) xor (layer2_outputs(636)));
    outputs(6122) <= not((layer2_outputs(2602)) xor (layer2_outputs(2978)));
    outputs(6123) <= layer2_outputs(4731);
    outputs(6124) <= not((layer2_outputs(2971)) and (layer2_outputs(5868)));
    outputs(6125) <= (layer2_outputs(7251)) xor (layer2_outputs(5187));
    outputs(6126) <= not(layer2_outputs(5645));
    outputs(6127) <= layer2_outputs(3996);
    outputs(6128) <= not(layer2_outputs(4003));
    outputs(6129) <= not((layer2_outputs(9701)) xor (layer2_outputs(7580)));
    outputs(6130) <= not((layer2_outputs(8675)) or (layer2_outputs(1718)));
    outputs(6131) <= not(layer2_outputs(9556));
    outputs(6132) <= layer2_outputs(7682);
    outputs(6133) <= not(layer2_outputs(2251));
    outputs(6134) <= (layer2_outputs(5032)) xor (layer2_outputs(6791));
    outputs(6135) <= not((layer2_outputs(5026)) xor (layer2_outputs(2857)));
    outputs(6136) <= layer2_outputs(2761);
    outputs(6137) <= (layer2_outputs(6656)) xor (layer2_outputs(9678));
    outputs(6138) <= not(layer2_outputs(3954));
    outputs(6139) <= layer2_outputs(2574);
    outputs(6140) <= not(layer2_outputs(7573));
    outputs(6141) <= not(layer2_outputs(3916));
    outputs(6142) <= not((layer2_outputs(3564)) xor (layer2_outputs(8044)));
    outputs(6143) <= not(layer2_outputs(10151));
    outputs(6144) <= layer2_outputs(5238);
    outputs(6145) <= not(layer2_outputs(4967));
    outputs(6146) <= not(layer2_outputs(10186));
    outputs(6147) <= layer2_outputs(3856);
    outputs(6148) <= (layer2_outputs(8447)) xor (layer2_outputs(3541));
    outputs(6149) <= not(layer2_outputs(2643));
    outputs(6150) <= not(layer2_outputs(339));
    outputs(6151) <= not(layer2_outputs(4332));
    outputs(6152) <= layer2_outputs(3044);
    outputs(6153) <= (layer2_outputs(4224)) and (layer2_outputs(7615));
    outputs(6154) <= layer2_outputs(7110);
    outputs(6155) <= layer2_outputs(5771);
    outputs(6156) <= (layer2_outputs(5558)) xor (layer2_outputs(2655));
    outputs(6157) <= (layer2_outputs(9723)) and not (layer2_outputs(4832));
    outputs(6158) <= (layer2_outputs(847)) xor (layer2_outputs(5985));
    outputs(6159) <= not((layer2_outputs(1618)) or (layer2_outputs(4437)));
    outputs(6160) <= not(layer2_outputs(1838));
    outputs(6161) <= layer2_outputs(2263);
    outputs(6162) <= layer2_outputs(2543);
    outputs(6163) <= not(layer2_outputs(6110));
    outputs(6164) <= not((layer2_outputs(382)) xor (layer2_outputs(2566)));
    outputs(6165) <= (layer2_outputs(9005)) and not (layer2_outputs(966));
    outputs(6166) <= not(layer2_outputs(784));
    outputs(6167) <= not(layer2_outputs(5192)) or (layer2_outputs(4431));
    outputs(6168) <= layer2_outputs(9671);
    outputs(6169) <= not((layer2_outputs(9123)) and (layer2_outputs(7917)));
    outputs(6170) <= not((layer2_outputs(8031)) and (layer2_outputs(6047)));
    outputs(6171) <= not(layer2_outputs(9144));
    outputs(6172) <= layer2_outputs(3799);
    outputs(6173) <= layer2_outputs(2695);
    outputs(6174) <= layer2_outputs(7076);
    outputs(6175) <= layer2_outputs(5442);
    outputs(6176) <= not(layer2_outputs(6351));
    outputs(6177) <= layer2_outputs(10165);
    outputs(6178) <= not(layer2_outputs(3228));
    outputs(6179) <= layer2_outputs(3722);
    outputs(6180) <= layer2_outputs(10191);
    outputs(6181) <= not(layer2_outputs(606));
    outputs(6182) <= not(layer2_outputs(3769));
    outputs(6183) <= not(layer2_outputs(4196));
    outputs(6184) <= not(layer2_outputs(9692));
    outputs(6185) <= not(layer2_outputs(6106));
    outputs(6186) <= not((layer2_outputs(6374)) xor (layer2_outputs(654)));
    outputs(6187) <= layer2_outputs(8003);
    outputs(6188) <= layer2_outputs(1736);
    outputs(6189) <= layer2_outputs(8274);
    outputs(6190) <= (layer2_outputs(4694)) xor (layer2_outputs(5769));
    outputs(6191) <= (layer2_outputs(6615)) and not (layer2_outputs(7312));
    outputs(6192) <= not(layer2_outputs(9644));
    outputs(6193) <= layer2_outputs(786);
    outputs(6194) <= not(layer2_outputs(9817));
    outputs(6195) <= (layer2_outputs(5314)) and not (layer2_outputs(2238));
    outputs(6196) <= (layer2_outputs(4134)) and (layer2_outputs(6001));
    outputs(6197) <= not(layer2_outputs(5676));
    outputs(6198) <= not(layer2_outputs(735));
    outputs(6199) <= not(layer2_outputs(6687));
    outputs(6200) <= (layer2_outputs(4925)) xor (layer2_outputs(7233));
    outputs(6201) <= not(layer2_outputs(1509));
    outputs(6202) <= not(layer2_outputs(5198));
    outputs(6203) <= not(layer2_outputs(8599));
    outputs(6204) <= not((layer2_outputs(4522)) xor (layer2_outputs(9472)));
    outputs(6205) <= (layer2_outputs(5426)) xor (layer2_outputs(6490));
    outputs(6206) <= not(layer2_outputs(9965));
    outputs(6207) <= not(layer2_outputs(360));
    outputs(6208) <= (layer2_outputs(9510)) xor (layer2_outputs(5463));
    outputs(6209) <= (layer2_outputs(1007)) and not (layer2_outputs(1695));
    outputs(6210) <= not((layer2_outputs(2892)) xor (layer2_outputs(8562)));
    outputs(6211) <= not((layer2_outputs(1235)) xor (layer2_outputs(7389)));
    outputs(6212) <= layer2_outputs(9210);
    outputs(6213) <= (layer2_outputs(9357)) xor (layer2_outputs(8419));
    outputs(6214) <= not((layer2_outputs(5875)) or (layer2_outputs(2035)));
    outputs(6215) <= not(layer2_outputs(8174));
    outputs(6216) <= layer2_outputs(6150);
    outputs(6217) <= (layer2_outputs(8196)) xor (layer2_outputs(9775));
    outputs(6218) <= not(layer2_outputs(2931));
    outputs(6219) <= (layer2_outputs(7246)) xor (layer2_outputs(6255));
    outputs(6220) <= layer2_outputs(9455);
    outputs(6221) <= layer2_outputs(1009);
    outputs(6222) <= layer2_outputs(3914);
    outputs(6223) <= (layer2_outputs(10072)) and (layer2_outputs(1635));
    outputs(6224) <= not((layer2_outputs(8555)) xor (layer2_outputs(6797)));
    outputs(6225) <= not(layer2_outputs(9375));
    outputs(6226) <= not(layer2_outputs(671));
    outputs(6227) <= (layer2_outputs(1194)) xor (layer2_outputs(6386));
    outputs(6228) <= not(layer2_outputs(2406));
    outputs(6229) <= not(layer2_outputs(4966));
    outputs(6230) <= not(layer2_outputs(4511));
    outputs(6231) <= (layer2_outputs(3311)) xor (layer2_outputs(6779));
    outputs(6232) <= layer2_outputs(1355);
    outputs(6233) <= not(layer2_outputs(8587));
    outputs(6234) <= not((layer2_outputs(5967)) xor (layer2_outputs(62)));
    outputs(6235) <= not((layer2_outputs(7480)) or (layer2_outputs(3954)));
    outputs(6236) <= layer2_outputs(4771);
    outputs(6237) <= not(layer2_outputs(1777));
    outputs(6238) <= layer2_outputs(7175);
    outputs(6239) <= (layer2_outputs(2599)) and not (layer2_outputs(1195));
    outputs(6240) <= layer2_outputs(8650);
    outputs(6241) <= not(layer2_outputs(6016));
    outputs(6242) <= layer2_outputs(2474);
    outputs(6243) <= (layer2_outputs(2312)) xor (layer2_outputs(7723));
    outputs(6244) <= (layer2_outputs(9934)) xor (layer2_outputs(2640));
    outputs(6245) <= not(layer2_outputs(7132));
    outputs(6246) <= not(layer2_outputs(3743));
    outputs(6247) <= layer2_outputs(9524);
    outputs(6248) <= not(layer2_outputs(8206));
    outputs(6249) <= layer2_outputs(2431);
    outputs(6250) <= (layer2_outputs(1467)) and (layer2_outputs(6812));
    outputs(6251) <= not((layer2_outputs(5597)) xor (layer2_outputs(8638)));
    outputs(6252) <= layer2_outputs(3847);
    outputs(6253) <= not(layer2_outputs(9623));
    outputs(6254) <= not(layer2_outputs(8303));
    outputs(6255) <= not(layer2_outputs(7122));
    outputs(6256) <= not(layer2_outputs(4157));
    outputs(6257) <= not((layer2_outputs(9538)) xor (layer2_outputs(52)));
    outputs(6258) <= not(layer2_outputs(7903));
    outputs(6259) <= layer2_outputs(1244);
    outputs(6260) <= (layer2_outputs(2631)) xor (layer2_outputs(5454));
    outputs(6261) <= not(layer2_outputs(4297));
    outputs(6262) <= (layer2_outputs(8027)) xor (layer2_outputs(10110));
    outputs(6263) <= layer2_outputs(5902);
    outputs(6264) <= layer2_outputs(7382);
    outputs(6265) <= (layer2_outputs(8637)) and not (layer2_outputs(7044));
    outputs(6266) <= not(layer2_outputs(7539));
    outputs(6267) <= not(layer2_outputs(6594));
    outputs(6268) <= layer2_outputs(9047);
    outputs(6269) <= not(layer2_outputs(6045));
    outputs(6270) <= not((layer2_outputs(4412)) xor (layer2_outputs(4600)));
    outputs(6271) <= not(layer2_outputs(300));
    outputs(6272) <= not((layer2_outputs(6650)) xor (layer2_outputs(7915)));
    outputs(6273) <= layer2_outputs(4928);
    outputs(6274) <= not(layer2_outputs(5880));
    outputs(6275) <= layer2_outputs(1418);
    outputs(6276) <= not(layer2_outputs(8222));
    outputs(6277) <= layer2_outputs(7481);
    outputs(6278) <= not((layer2_outputs(6690)) xor (layer2_outputs(6084)));
    outputs(6279) <= (layer2_outputs(5027)) xor (layer2_outputs(7339));
    outputs(6280) <= layer2_outputs(5118);
    outputs(6281) <= not(layer2_outputs(239));
    outputs(6282) <= not(layer2_outputs(1792));
    outputs(6283) <= (layer2_outputs(2492)) and not (layer2_outputs(7609));
    outputs(6284) <= not((layer2_outputs(8173)) xor (layer2_outputs(7871)));
    outputs(6285) <= layer2_outputs(1939);
    outputs(6286) <= layer2_outputs(6215);
    outputs(6287) <= layer2_outputs(959);
    outputs(6288) <= not(layer2_outputs(4765));
    outputs(6289) <= not((layer2_outputs(7233)) xor (layer2_outputs(2413)));
    outputs(6290) <= (layer2_outputs(6414)) xor (layer2_outputs(4189));
    outputs(6291) <= (layer2_outputs(9370)) xor (layer2_outputs(1664));
    outputs(6292) <= not((layer2_outputs(871)) xor (layer2_outputs(3362)));
    outputs(6293) <= not(layer2_outputs(6548));
    outputs(6294) <= layer2_outputs(4167);
    outputs(6295) <= not(layer2_outputs(1310));
    outputs(6296) <= not(layer2_outputs(8574));
    outputs(6297) <= layer2_outputs(8592);
    outputs(6298) <= not(layer2_outputs(9227));
    outputs(6299) <= not(layer2_outputs(9566));
    outputs(6300) <= not((layer2_outputs(5153)) xor (layer2_outputs(7654)));
    outputs(6301) <= not(layer2_outputs(4143));
    outputs(6302) <= (layer2_outputs(4299)) and not (layer2_outputs(10202));
    outputs(6303) <= not((layer2_outputs(5761)) xor (layer2_outputs(8774)));
    outputs(6304) <= not((layer2_outputs(9319)) xor (layer2_outputs(2601)));
    outputs(6305) <= (layer2_outputs(982)) xor (layer2_outputs(8833));
    outputs(6306) <= not((layer2_outputs(9937)) xor (layer2_outputs(2979)));
    outputs(6307) <= (layer2_outputs(878)) and (layer2_outputs(2891));
    outputs(6308) <= not((layer2_outputs(1079)) xor (layer2_outputs(1178)));
    outputs(6309) <= (layer2_outputs(3305)) and (layer2_outputs(8673));
    outputs(6310) <= (layer2_outputs(7121)) and not (layer2_outputs(4911));
    outputs(6311) <= layer2_outputs(8780);
    outputs(6312) <= layer2_outputs(2569);
    outputs(6313) <= not(layer2_outputs(7831));
    outputs(6314) <= (layer2_outputs(3173)) and not (layer2_outputs(7502));
    outputs(6315) <= layer2_outputs(5342);
    outputs(6316) <= layer2_outputs(7764);
    outputs(6317) <= layer2_outputs(9581);
    outputs(6318) <= layer2_outputs(9521);
    outputs(6319) <= not(layer2_outputs(8972));
    outputs(6320) <= (layer2_outputs(9239)) xor (layer2_outputs(1167));
    outputs(6321) <= not(layer2_outputs(9376)) or (layer2_outputs(4104));
    outputs(6322) <= layer2_outputs(7425);
    outputs(6323) <= (layer2_outputs(7999)) and not (layer2_outputs(8500));
    outputs(6324) <= layer2_outputs(6223);
    outputs(6325) <= layer2_outputs(10117);
    outputs(6326) <= not(layer2_outputs(3063));
    outputs(6327) <= layer2_outputs(7418);
    outputs(6328) <= layer2_outputs(8920);
    outputs(6329) <= not(layer2_outputs(1050));
    outputs(6330) <= not((layer2_outputs(9724)) xor (layer2_outputs(10215)));
    outputs(6331) <= not(layer2_outputs(9175));
    outputs(6332) <= layer2_outputs(8586);
    outputs(6333) <= not((layer2_outputs(7348)) and (layer2_outputs(10176)));
    outputs(6334) <= layer2_outputs(10128);
    outputs(6335) <= layer2_outputs(7621);
    outputs(6336) <= layer2_outputs(7116);
    outputs(6337) <= layer2_outputs(8199);
    outputs(6338) <= not(layer2_outputs(8705)) or (layer2_outputs(6355));
    outputs(6339) <= layer2_outputs(2184);
    outputs(6340) <= layer2_outputs(8336);
    outputs(6341) <= (layer2_outputs(429)) and not (layer2_outputs(3938));
    outputs(6342) <= not(layer2_outputs(1618));
    outputs(6343) <= not(layer2_outputs(7592));
    outputs(6344) <= not(layer2_outputs(7006));
    outputs(6345) <= (layer2_outputs(9408)) and not (layer2_outputs(551));
    outputs(6346) <= (layer2_outputs(2145)) xor (layer2_outputs(864));
    outputs(6347) <= layer2_outputs(7113);
    outputs(6348) <= not(layer2_outputs(6935));
    outputs(6349) <= not(layer2_outputs(5484));
    outputs(6350) <= not(layer2_outputs(9635));
    outputs(6351) <= layer2_outputs(6019);
    outputs(6352) <= not(layer2_outputs(1528));
    outputs(6353) <= layer2_outputs(6942);
    outputs(6354) <= not(layer2_outputs(4314)) or (layer2_outputs(4703));
    outputs(6355) <= not((layer2_outputs(7071)) or (layer2_outputs(3888)));
    outputs(6356) <= layer2_outputs(1531);
    outputs(6357) <= (layer2_outputs(8613)) and not (layer2_outputs(8417));
    outputs(6358) <= not((layer2_outputs(3718)) xor (layer2_outputs(4036)));
    outputs(6359) <= not(layer2_outputs(1970));
    outputs(6360) <= (layer2_outputs(6105)) xor (layer2_outputs(5044));
    outputs(6361) <= not((layer2_outputs(5220)) or (layer2_outputs(7800)));
    outputs(6362) <= layer2_outputs(9772);
    outputs(6363) <= layer2_outputs(9976);
    outputs(6364) <= (layer2_outputs(6819)) and not (layer2_outputs(5439));
    outputs(6365) <= not(layer2_outputs(7061));
    outputs(6366) <= not(layer2_outputs(954));
    outputs(6367) <= not((layer2_outputs(6424)) xor (layer2_outputs(8438)));
    outputs(6368) <= layer2_outputs(9358);
    outputs(6369) <= layer2_outputs(812);
    outputs(6370) <= layer2_outputs(8110);
    outputs(6371) <= not(layer2_outputs(9939));
    outputs(6372) <= (layer2_outputs(164)) xor (layer2_outputs(1408));
    outputs(6373) <= not(layer2_outputs(3257));
    outputs(6374) <= layer2_outputs(35);
    outputs(6375) <= (layer2_outputs(4673)) xor (layer2_outputs(8417));
    outputs(6376) <= not(layer2_outputs(1845));
    outputs(6377) <= not(layer2_outputs(971)) or (layer2_outputs(3326));
    outputs(6378) <= not(layer2_outputs(2344));
    outputs(6379) <= not(layer2_outputs(507));
    outputs(6380) <= not(layer2_outputs(1623));
    outputs(6381) <= (layer2_outputs(5811)) and not (layer2_outputs(5230));
    outputs(6382) <= layer2_outputs(6079);
    outputs(6383) <= not(layer2_outputs(3019));
    outputs(6384) <= not(layer2_outputs(3052)) or (layer2_outputs(637));
    outputs(6385) <= layer2_outputs(2020);
    outputs(6386) <= not(layer2_outputs(8532));
    outputs(6387) <= not(layer2_outputs(7457));
    outputs(6388) <= (layer2_outputs(1677)) xor (layer2_outputs(5997));
    outputs(6389) <= not(layer2_outputs(4188));
    outputs(6390) <= not(layer2_outputs(8451));
    outputs(6391) <= (layer2_outputs(223)) xor (layer2_outputs(6723));
    outputs(6392) <= (layer2_outputs(9756)) xor (layer2_outputs(694));
    outputs(6393) <= not(layer2_outputs(4870));
    outputs(6394) <= layer2_outputs(5410);
    outputs(6395) <= not(layer2_outputs(6387));
    outputs(6396) <= not(layer2_outputs(3882));
    outputs(6397) <= (layer2_outputs(8775)) xor (layer2_outputs(9512));
    outputs(6398) <= (layer2_outputs(4815)) and (layer2_outputs(3999));
    outputs(6399) <= (layer2_outputs(3226)) and not (layer2_outputs(5047));
    outputs(6400) <= not(layer2_outputs(971));
    outputs(6401) <= layer2_outputs(3318);
    outputs(6402) <= not((layer2_outputs(9231)) xor (layer2_outputs(1572)));
    outputs(6403) <= not(layer2_outputs(4835));
    outputs(6404) <= not((layer2_outputs(3145)) or (layer2_outputs(1502)));
    outputs(6405) <= layer2_outputs(6191);
    outputs(6406) <= (layer2_outputs(6749)) or (layer2_outputs(6677));
    outputs(6407) <= layer2_outputs(7684);
    outputs(6408) <= not(layer2_outputs(8721));
    outputs(6409) <= layer2_outputs(1137);
    outputs(6410) <= not(layer2_outputs(4579)) or (layer2_outputs(9987));
    outputs(6411) <= layer2_outputs(1712);
    outputs(6412) <= not((layer2_outputs(4310)) xor (layer2_outputs(6508)));
    outputs(6413) <= not((layer2_outputs(6403)) or (layer2_outputs(8356)));
    outputs(6414) <= not(layer2_outputs(8396));
    outputs(6415) <= not((layer2_outputs(1096)) xor (layer2_outputs(6997)));
    outputs(6416) <= (layer2_outputs(7446)) or (layer2_outputs(4797));
    outputs(6417) <= not(layer2_outputs(5155));
    outputs(6418) <= layer2_outputs(1873);
    outputs(6419) <= not((layer2_outputs(2854)) or (layer2_outputs(5765)));
    outputs(6420) <= layer2_outputs(1145);
    outputs(6421) <= not(layer2_outputs(6232));
    outputs(6422) <= not(layer2_outputs(5805)) or (layer2_outputs(8845));
    outputs(6423) <= not(layer2_outputs(1648));
    outputs(6424) <= (layer2_outputs(5333)) and not (layer2_outputs(2693));
    outputs(6425) <= not((layer2_outputs(9569)) or (layer2_outputs(129)));
    outputs(6426) <= layer2_outputs(7861);
    outputs(6427) <= not(layer2_outputs(8426));
    outputs(6428) <= (layer2_outputs(5536)) xor (layer2_outputs(2367));
    outputs(6429) <= not(layer2_outputs(4728)) or (layer2_outputs(7405));
    outputs(6430) <= layer2_outputs(9520);
    outputs(6431) <= not((layer2_outputs(9263)) or (layer2_outputs(8546)));
    outputs(6432) <= not(layer2_outputs(9862)) or (layer2_outputs(1057));
    outputs(6433) <= not(layer2_outputs(2546));
    outputs(6434) <= layer2_outputs(2820);
    outputs(6435) <= not(layer2_outputs(2522));
    outputs(6436) <= not(layer2_outputs(1727));
    outputs(6437) <= not(layer2_outputs(4205));
    outputs(6438) <= not((layer2_outputs(4686)) xor (layer2_outputs(5223)));
    outputs(6439) <= not(layer2_outputs(5129));
    outputs(6440) <= not(layer2_outputs(9755));
    outputs(6441) <= not(layer2_outputs(9843));
    outputs(6442) <= layer2_outputs(9022);
    outputs(6443) <= layer2_outputs(5591);
    outputs(6444) <= not((layer2_outputs(8743)) xor (layer2_outputs(3916)));
    outputs(6445) <= not((layer2_outputs(3089)) or (layer2_outputs(5334)));
    outputs(6446) <= layer2_outputs(6550);
    outputs(6447) <= (layer2_outputs(6640)) xor (layer2_outputs(4132));
    outputs(6448) <= layer2_outputs(5149);
    outputs(6449) <= not(layer2_outputs(8215));
    outputs(6450) <= not((layer2_outputs(7548)) xor (layer2_outputs(4122)));
    outputs(6451) <= layer2_outputs(9447);
    outputs(6452) <= not(layer2_outputs(9343));
    outputs(6453) <= (layer2_outputs(5843)) and not (layer2_outputs(3510));
    outputs(6454) <= layer2_outputs(5538);
    outputs(6455) <= (layer2_outputs(7575)) and (layer2_outputs(9359));
    outputs(6456) <= layer2_outputs(2073);
    outputs(6457) <= (layer2_outputs(1843)) and not (layer2_outputs(338));
    outputs(6458) <= not(layer2_outputs(874));
    outputs(6459) <= (layer2_outputs(4653)) and not (layer2_outputs(4892));
    outputs(6460) <= not(layer2_outputs(581));
    outputs(6461) <= not(layer2_outputs(6738));
    outputs(6462) <= not(layer2_outputs(3400));
    outputs(6463) <= (layer2_outputs(38)) or (layer2_outputs(2012));
    outputs(6464) <= layer2_outputs(894);
    outputs(6465) <= layer2_outputs(6668);
    outputs(6466) <= (layer2_outputs(3174)) and (layer2_outputs(4350));
    outputs(6467) <= not(layer2_outputs(6941));
    outputs(6468) <= not((layer2_outputs(2984)) xor (layer2_outputs(6072)));
    outputs(6469) <= not(layer2_outputs(4940));
    outputs(6470) <= not(layer2_outputs(8905));
    outputs(6471) <= not(layer2_outputs(362));
    outputs(6472) <= not((layer2_outputs(7048)) or (layer2_outputs(6970)));
    outputs(6473) <= (layer2_outputs(9453)) and not (layer2_outputs(8312));
    outputs(6474) <= layer2_outputs(1646);
    outputs(6475) <= layer2_outputs(226);
    outputs(6476) <= not(layer2_outputs(2089));
    outputs(6477) <= not((layer2_outputs(1149)) or (layer2_outputs(1469)));
    outputs(6478) <= (layer2_outputs(1602)) and not (layer2_outputs(7398));
    outputs(6479) <= not((layer2_outputs(3350)) xor (layer2_outputs(3075)));
    outputs(6480) <= layer2_outputs(6829);
    outputs(6481) <= layer2_outputs(1282);
    outputs(6482) <= layer2_outputs(6003);
    outputs(6483) <= (layer2_outputs(1593)) xor (layer2_outputs(2757));
    outputs(6484) <= not(layer2_outputs(7635));
    outputs(6485) <= not(layer2_outputs(9782));
    outputs(6486) <= not((layer2_outputs(6616)) xor (layer2_outputs(2647)));
    outputs(6487) <= not(layer2_outputs(4663));
    outputs(6488) <= not((layer2_outputs(466)) xor (layer2_outputs(9978)));
    outputs(6489) <= (layer2_outputs(5409)) and not (layer2_outputs(8925));
    outputs(6490) <= not(layer2_outputs(8853));
    outputs(6491) <= layer2_outputs(2206);
    outputs(6492) <= (layer2_outputs(3887)) and not (layer2_outputs(2789));
    outputs(6493) <= not(layer2_outputs(1767));
    outputs(6494) <= layer2_outputs(3958);
    outputs(6495) <= layer2_outputs(9048);
    outputs(6496) <= not(layer2_outputs(4128));
    outputs(6497) <= not(layer2_outputs(9331)) or (layer2_outputs(5617));
    outputs(6498) <= (layer2_outputs(1279)) xor (layer2_outputs(9636));
    outputs(6499) <= not((layer2_outputs(8684)) xor (layer2_outputs(7210)));
    outputs(6500) <= layer2_outputs(2086);
    outputs(6501) <= not(layer2_outputs(7631));
    outputs(6502) <= layer2_outputs(5816);
    outputs(6503) <= layer2_outputs(4981);
    outputs(6504) <= not((layer2_outputs(10051)) xor (layer2_outputs(1800)));
    outputs(6505) <= layer2_outputs(3610);
    outputs(6506) <= not((layer2_outputs(1989)) and (layer2_outputs(3754)));
    outputs(6507) <= not(layer2_outputs(6750));
    outputs(6508) <= not(layer2_outputs(5478));
    outputs(6509) <= layer2_outputs(10226);
    outputs(6510) <= layer2_outputs(8277);
    outputs(6511) <= not(layer2_outputs(10010));
    outputs(6512) <= not(layer2_outputs(9763));
    outputs(6513) <= layer2_outputs(6217);
    outputs(6514) <= not(layer2_outputs(4187));
    outputs(6515) <= not(layer2_outputs(5481));
    outputs(6516) <= not((layer2_outputs(8685)) xor (layer2_outputs(1620)));
    outputs(6517) <= layer2_outputs(7476);
    outputs(6518) <= not(layer2_outputs(6469));
    outputs(6519) <= layer2_outputs(4901);
    outputs(6520) <= not(layer2_outputs(6859));
    outputs(6521) <= not(layer2_outputs(4153));
    outputs(6522) <= not(layer2_outputs(9102));
    outputs(6523) <= layer2_outputs(6192);
    outputs(6524) <= (layer2_outputs(6547)) and (layer2_outputs(4149));
    outputs(6525) <= layer2_outputs(4877);
    outputs(6526) <= layer2_outputs(5648);
    outputs(6527) <= not(layer2_outputs(7719));
    outputs(6528) <= not(layer2_outputs(2015));
    outputs(6529) <= layer2_outputs(1839);
    outputs(6530) <= not(layer2_outputs(9691));
    outputs(6531) <= not((layer2_outputs(2583)) xor (layer2_outputs(8542)));
    outputs(6532) <= not(layer2_outputs(8466));
    outputs(6533) <= layer2_outputs(3666);
    outputs(6534) <= layer2_outputs(8918);
    outputs(6535) <= not((layer2_outputs(5434)) xor (layer2_outputs(9253)));
    outputs(6536) <= not((layer2_outputs(6979)) and (layer2_outputs(10210)));
    outputs(6537) <= not(layer2_outputs(1648));
    outputs(6538) <= layer2_outputs(264);
    outputs(6539) <= not(layer2_outputs(5966));
    outputs(6540) <= not(layer2_outputs(3694));
    outputs(6541) <= not((layer2_outputs(9135)) and (layer2_outputs(3649)));
    outputs(6542) <= layer2_outputs(471);
    outputs(6543) <= (layer2_outputs(3737)) and not (layer2_outputs(3623));
    outputs(6544) <= layer2_outputs(7095);
    outputs(6545) <= layer2_outputs(6864);
    outputs(6546) <= (layer2_outputs(4474)) and (layer2_outputs(5269));
    outputs(6547) <= layer2_outputs(2208);
    outputs(6548) <= not(layer2_outputs(8178));
    outputs(6549) <= (layer2_outputs(5439)) xor (layer2_outputs(8374));
    outputs(6550) <= not(layer2_outputs(2080));
    outputs(6551) <= not((layer2_outputs(3630)) or (layer2_outputs(5750)));
    outputs(6552) <= layer2_outputs(6628);
    outputs(6553) <= (layer2_outputs(6988)) and not (layer2_outputs(8722));
    outputs(6554) <= layer2_outputs(9434);
    outputs(6555) <= not((layer2_outputs(1431)) or (layer2_outputs(8897)));
    outputs(6556) <= layer2_outputs(2945);
    outputs(6557) <= not((layer2_outputs(6185)) xor (layer2_outputs(4413)));
    outputs(6558) <= layer2_outputs(9399);
    outputs(6559) <= (layer2_outputs(4772)) xor (layer2_outputs(4075));
    outputs(6560) <= layer2_outputs(1457);
    outputs(6561) <= layer2_outputs(2777);
    outputs(6562) <= not(layer2_outputs(152));
    outputs(6563) <= not(layer2_outputs(7763));
    outputs(6564) <= layer2_outputs(1063);
    outputs(6565) <= not((layer2_outputs(9598)) or (layer2_outputs(347)));
    outputs(6566) <= not(layer2_outputs(1852));
    outputs(6567) <= not(layer2_outputs(8949));
    outputs(6568) <= layer2_outputs(4215);
    outputs(6569) <= not(layer2_outputs(8256));
    outputs(6570) <= layer2_outputs(4711);
    outputs(6571) <= layer2_outputs(717);
    outputs(6572) <= layer2_outputs(2379);
    outputs(6573) <= not(layer2_outputs(9653));
    outputs(6574) <= not(layer2_outputs(322));
    outputs(6575) <= layer2_outputs(3565);
    outputs(6576) <= (layer2_outputs(6122)) xor (layer2_outputs(3811));
    outputs(6577) <= (layer2_outputs(3501)) xor (layer2_outputs(4697));
    outputs(6578) <= layer2_outputs(3955);
    outputs(6579) <= (layer2_outputs(2794)) or (layer2_outputs(3279));
    outputs(6580) <= not(layer2_outputs(1186)) or (layer2_outputs(1526));
    outputs(6581) <= not(layer2_outputs(1727));
    outputs(6582) <= not(layer2_outputs(9464));
    outputs(6583) <= (layer2_outputs(1008)) or (layer2_outputs(156));
    outputs(6584) <= (layer2_outputs(2217)) or (layer2_outputs(8520));
    outputs(6585) <= not((layer2_outputs(6410)) xor (layer2_outputs(1738)));
    outputs(6586) <= layer2_outputs(790);
    outputs(6587) <= not(layer2_outputs(7671)) or (layer2_outputs(5749));
    outputs(6588) <= layer2_outputs(6008);
    outputs(6589) <= not(layer2_outputs(6059));
    outputs(6590) <= layer2_outputs(9401);
    outputs(6591) <= layer2_outputs(5388);
    outputs(6592) <= (layer2_outputs(9161)) xor (layer2_outputs(902));
    outputs(6593) <= not((layer2_outputs(6696)) or (layer2_outputs(8047)));
    outputs(6594) <= not(layer2_outputs(1026));
    outputs(6595) <= not(layer2_outputs(2368));
    outputs(6596) <= layer2_outputs(5097);
    outputs(6597) <= layer2_outputs(1540);
    outputs(6598) <= layer2_outputs(8651);
    outputs(6599) <= not((layer2_outputs(6088)) or (layer2_outputs(4568)));
    outputs(6600) <= not((layer2_outputs(8683)) xor (layer2_outputs(2826)));
    outputs(6601) <= not(layer2_outputs(7984));
    outputs(6602) <= not((layer2_outputs(7746)) xor (layer2_outputs(4702)));
    outputs(6603) <= (layer2_outputs(8519)) and not (layer2_outputs(3706));
    outputs(6604) <= not((layer2_outputs(4488)) xor (layer2_outputs(8210)));
    outputs(6605) <= (layer2_outputs(8741)) xor (layer2_outputs(4432));
    outputs(6606) <= layer2_outputs(3210);
    outputs(6607) <= not(layer2_outputs(9405));
    outputs(6608) <= not((layer2_outputs(8243)) and (layer2_outputs(173)));
    outputs(6609) <= (layer2_outputs(5988)) and (layer2_outputs(9724));
    outputs(6610) <= not((layer2_outputs(7473)) or (layer2_outputs(3476)));
    outputs(6611) <= not((layer2_outputs(2556)) xor (layer2_outputs(8192)));
    outputs(6612) <= layer2_outputs(1094);
    outputs(6613) <= not(layer2_outputs(7895));
    outputs(6614) <= (layer2_outputs(764)) or (layer2_outputs(8049));
    outputs(6615) <= layer2_outputs(9388);
    outputs(6616) <= not(layer2_outputs(5228));
    outputs(6617) <= layer2_outputs(103);
    outputs(6618) <= not(layer2_outputs(6722)) or (layer2_outputs(3188));
    outputs(6619) <= not(layer2_outputs(6888));
    outputs(6620) <= layer2_outputs(4904);
    outputs(6621) <= not((layer2_outputs(6509)) xor (layer2_outputs(7383)));
    outputs(6622) <= not(layer2_outputs(2164));
    outputs(6623) <= not((layer2_outputs(104)) xor (layer2_outputs(3763)));
    outputs(6624) <= not(layer2_outputs(8045));
    outputs(6625) <= layer2_outputs(6624);
    outputs(6626) <= layer2_outputs(6095);
    outputs(6627) <= not((layer2_outputs(1595)) xor (layer2_outputs(465)));
    outputs(6628) <= layer2_outputs(9942);
    outputs(6629) <= layer2_outputs(2541);
    outputs(6630) <= not(layer2_outputs(4102));
    outputs(6631) <= not(layer2_outputs(2450));
    outputs(6632) <= layer2_outputs(9707);
    outputs(6633) <= not(layer2_outputs(2518)) or (layer2_outputs(844));
    outputs(6634) <= (layer2_outputs(8084)) xor (layer2_outputs(7920));
    outputs(6635) <= not(layer2_outputs(2782));
    outputs(6636) <= layer2_outputs(2703);
    outputs(6637) <= (layer2_outputs(4653)) and not (layer2_outputs(614));
    outputs(6638) <= layer2_outputs(9301);
    outputs(6639) <= not((layer2_outputs(4896)) xor (layer2_outputs(1854)));
    outputs(6640) <= layer2_outputs(3551);
    outputs(6641) <= layer2_outputs(6621);
    outputs(6642) <= layer2_outputs(7544);
    outputs(6643) <= not(layer2_outputs(7842));
    outputs(6644) <= layer2_outputs(5623);
    outputs(6645) <= not((layer2_outputs(2036)) or (layer2_outputs(1376)));
    outputs(6646) <= layer2_outputs(5892);
    outputs(6647) <= layer2_outputs(6524);
    outputs(6648) <= not(layer2_outputs(597));
    outputs(6649) <= layer2_outputs(8487);
    outputs(6650) <= layer2_outputs(5716);
    outputs(6651) <= not(layer2_outputs(574));
    outputs(6652) <= not(layer2_outputs(9858));
    outputs(6653) <= not(layer2_outputs(5018));
    outputs(6654) <= layer2_outputs(9434);
    outputs(6655) <= not(layer2_outputs(9924));
    outputs(6656) <= not(layer2_outputs(2007));
    outputs(6657) <= not(layer2_outputs(3032));
    outputs(6658) <= layer2_outputs(1652);
    outputs(6659) <= (layer2_outputs(8801)) and not (layer2_outputs(5501));
    outputs(6660) <= not(layer2_outputs(8500));
    outputs(6661) <= layer2_outputs(452);
    outputs(6662) <= not(layer2_outputs(7559)) or (layer2_outputs(1535));
    outputs(6663) <= not((layer2_outputs(2499)) xor (layer2_outputs(8132)));
    outputs(6664) <= not(layer2_outputs(5150));
    outputs(6665) <= (layer2_outputs(6849)) xor (layer2_outputs(2637));
    outputs(6666) <= (layer2_outputs(9758)) xor (layer2_outputs(2069));
    outputs(6667) <= not(layer2_outputs(6117));
    outputs(6668) <= (layer2_outputs(2186)) xor (layer2_outputs(716));
    outputs(6669) <= layer2_outputs(2837);
    outputs(6670) <= (layer2_outputs(547)) and not (layer2_outputs(6475));
    outputs(6671) <= not(layer2_outputs(8942));
    outputs(6672) <= layer2_outputs(4260);
    outputs(6673) <= layer2_outputs(8236);
    outputs(6674) <= layer2_outputs(8811);
    outputs(6675) <= not(layer2_outputs(106));
    outputs(6676) <= layer2_outputs(7415);
    outputs(6677) <= not((layer2_outputs(7558)) xor (layer2_outputs(9404)));
    outputs(6678) <= not(layer2_outputs(7530));
    outputs(6679) <= (layer2_outputs(1064)) xor (layer2_outputs(2125));
    outputs(6680) <= not(layer2_outputs(1216));
    outputs(6681) <= not(layer2_outputs(1777));
    outputs(6682) <= not(layer2_outputs(1924));
    outputs(6683) <= not(layer2_outputs(6567));
    outputs(6684) <= (layer2_outputs(5837)) and not (layer2_outputs(6714));
    outputs(6685) <= layer2_outputs(10102);
    outputs(6686) <= layer2_outputs(9559);
    outputs(6687) <= (layer2_outputs(7110)) xor (layer2_outputs(2058));
    outputs(6688) <= (layer2_outputs(5757)) and (layer2_outputs(8527));
    outputs(6689) <= not(layer2_outputs(1337));
    outputs(6690) <= layer2_outputs(6369);
    outputs(6691) <= layer2_outputs(9296);
    outputs(6692) <= not(layer2_outputs(9489));
    outputs(6693) <= (layer2_outputs(2470)) and not (layer2_outputs(25));
    outputs(6694) <= not(layer2_outputs(9004));
    outputs(6695) <= not(layer2_outputs(8502));
    outputs(6696) <= layer2_outputs(9513);
    outputs(6697) <= layer2_outputs(2897);
    outputs(6698) <= layer2_outputs(8217);
    outputs(6699) <= layer2_outputs(6352);
    outputs(6700) <= not((layer2_outputs(8191)) xor (layer2_outputs(8605)));
    outputs(6701) <= not(layer2_outputs(990));
    outputs(6702) <= layer2_outputs(7430);
    outputs(6703) <= layer2_outputs(3427);
    outputs(6704) <= not((layer2_outputs(4451)) xor (layer2_outputs(796)));
    outputs(6705) <= not((layer2_outputs(463)) xor (layer2_outputs(2188)));
    outputs(6706) <= not(layer2_outputs(2434));
    outputs(6707) <= not(layer2_outputs(5180));
    outputs(6708) <= (layer2_outputs(3424)) and not (layer2_outputs(7230));
    outputs(6709) <= (layer2_outputs(9220)) xor (layer2_outputs(7788));
    outputs(6710) <= not(layer2_outputs(8334));
    outputs(6711) <= layer2_outputs(7010);
    outputs(6712) <= not(layer2_outputs(10105));
    outputs(6713) <= (layer2_outputs(1612)) or (layer2_outputs(3651));
    outputs(6714) <= layer2_outputs(8348);
    outputs(6715) <= not(layer2_outputs(4463)) or (layer2_outputs(1120));
    outputs(6716) <= layer2_outputs(2437);
    outputs(6717) <= not(layer2_outputs(7250));
    outputs(6718) <= not(layer2_outputs(7050));
    outputs(6719) <= not((layer2_outputs(6609)) xor (layer2_outputs(9802)));
    outputs(6720) <= layer2_outputs(1700);
    outputs(6721) <= not((layer2_outputs(4495)) xor (layer2_outputs(2779)));
    outputs(6722) <= not(layer2_outputs(6070));
    outputs(6723) <= not(layer2_outputs(1755)) or (layer2_outputs(2135));
    outputs(6724) <= not((layer2_outputs(15)) xor (layer2_outputs(8400)));
    outputs(6725) <= layer2_outputs(9780);
    outputs(6726) <= (layer2_outputs(5918)) and (layer2_outputs(2063));
    outputs(6727) <= not((layer2_outputs(5678)) and (layer2_outputs(8574)));
    outputs(6728) <= not((layer2_outputs(16)) or (layer2_outputs(7970)));
    outputs(6729) <= not(layer2_outputs(7817));
    outputs(6730) <= layer2_outputs(7734);
    outputs(6731) <= not(layer2_outputs(2348));
    outputs(6732) <= layer2_outputs(4419);
    outputs(6733) <= not(layer2_outputs(7778));
    outputs(6734) <= not((layer2_outputs(3643)) xor (layer2_outputs(7231)));
    outputs(6735) <= (layer2_outputs(6422)) or (layer2_outputs(5149));
    outputs(6736) <= layer2_outputs(431);
    outputs(6737) <= not(layer2_outputs(2304));
    outputs(6738) <= not((layer2_outputs(6274)) xor (layer2_outputs(9000)));
    outputs(6739) <= not(layer2_outputs(6806));
    outputs(6740) <= layer2_outputs(6010);
    outputs(6741) <= not((layer2_outputs(182)) xor (layer2_outputs(8866)));
    outputs(6742) <= not(layer2_outputs(8181));
    outputs(6743) <= not(layer2_outputs(1404));
    outputs(6744) <= layer2_outputs(4465);
    outputs(6745) <= layer2_outputs(10171);
    outputs(6746) <= layer2_outputs(2735);
    outputs(6747) <= not((layer2_outputs(6475)) xor (layer2_outputs(5958)));
    outputs(6748) <= not(layer2_outputs(3727));
    outputs(6749) <= layer2_outputs(5360);
    outputs(6750) <= not(layer2_outputs(5629)) or (layer2_outputs(6462));
    outputs(6751) <= layer2_outputs(9402);
    outputs(6752) <= layer2_outputs(5904);
    outputs(6753) <= layer2_outputs(9916);
    outputs(6754) <= layer2_outputs(4595);
    outputs(6755) <= not(layer2_outputs(4897));
    outputs(6756) <= layer2_outputs(9596);
    outputs(6757) <= not(layer2_outputs(7839)) or (layer2_outputs(4345));
    outputs(6758) <= layer2_outputs(6452);
    outputs(6759) <= layer2_outputs(7879);
    outputs(6760) <= not(layer2_outputs(6432));
    outputs(6761) <= not(layer2_outputs(3190));
    outputs(6762) <= not(layer2_outputs(259));
    outputs(6763) <= not(layer2_outputs(2031));
    outputs(6764) <= layer2_outputs(3908);
    outputs(6765) <= layer2_outputs(353);
    outputs(6766) <= layer2_outputs(8939);
    outputs(6767) <= (layer2_outputs(42)) and not (layer2_outputs(7363));
    outputs(6768) <= not(layer2_outputs(575));
    outputs(6769) <= (layer2_outputs(3033)) xor (layer2_outputs(8615));
    outputs(6770) <= (layer2_outputs(346)) xor (layer2_outputs(2923));
    outputs(6771) <= layer2_outputs(3818);
    outputs(6772) <= not(layer2_outputs(10144));
    outputs(6773) <= layer2_outputs(125);
    outputs(6774) <= layer2_outputs(997);
    outputs(6775) <= layer2_outputs(7203);
    outputs(6776) <= layer2_outputs(2636);
    outputs(6777) <= not(layer2_outputs(2172)) or (layer2_outputs(3744));
    outputs(6778) <= (layer2_outputs(8449)) xor (layer2_outputs(9733));
    outputs(6779) <= not(layer2_outputs(9135)) or (layer2_outputs(3658));
    outputs(6780) <= (layer2_outputs(931)) or (layer2_outputs(624));
    outputs(6781) <= not(layer2_outputs(7745));
    outputs(6782) <= not(layer2_outputs(5933));
    outputs(6783) <= not((layer2_outputs(6571)) and (layer2_outputs(804)));
    outputs(6784) <= (layer2_outputs(8668)) xor (layer2_outputs(3019));
    outputs(6785) <= layer2_outputs(4401);
    outputs(6786) <= layer2_outputs(9438);
    outputs(6787) <= layer2_outputs(9415);
    outputs(6788) <= not(layer2_outputs(3219));
    outputs(6789) <= not(layer2_outputs(4503));
    outputs(6790) <= not(layer2_outputs(7417));
    outputs(6791) <= not(layer2_outputs(6104));
    outputs(6792) <= not((layer2_outputs(8041)) or (layer2_outputs(6255)));
    outputs(6793) <= layer2_outputs(166);
    outputs(6794) <= layer2_outputs(4923);
    outputs(6795) <= layer2_outputs(5443);
    outputs(6796) <= (layer2_outputs(6096)) and not (layer2_outputs(61));
    outputs(6797) <= layer2_outputs(8995);
    outputs(6798) <= layer2_outputs(2257);
    outputs(6799) <= (layer2_outputs(8379)) xor (layer2_outputs(3397));
    outputs(6800) <= (layer2_outputs(1312)) or (layer2_outputs(5499));
    outputs(6801) <= not(layer2_outputs(3292));
    outputs(6802) <= not((layer2_outputs(3740)) xor (layer2_outputs(3231)));
    outputs(6803) <= layer2_outputs(3087);
    outputs(6804) <= (layer2_outputs(5421)) xor (layer2_outputs(9248));
    outputs(6805) <= not(layer2_outputs(7138));
    outputs(6806) <= layer2_outputs(478);
    outputs(6807) <= layer2_outputs(5141);
    outputs(6808) <= not(layer2_outputs(3436));
    outputs(6809) <= not(layer2_outputs(6458)) or (layer2_outputs(2951));
    outputs(6810) <= (layer2_outputs(72)) and not (layer2_outputs(2736));
    outputs(6811) <= (layer2_outputs(7925)) xor (layer2_outputs(2937));
    outputs(6812) <= not(layer2_outputs(6197));
    outputs(6813) <= layer2_outputs(8398);
    outputs(6814) <= not((layer2_outputs(3825)) or (layer2_outputs(5219)));
    outputs(6815) <= (layer2_outputs(5959)) xor (layer2_outputs(8078));
    outputs(6816) <= (layer2_outputs(7035)) or (layer2_outputs(6652));
    outputs(6817) <= layer2_outputs(4385);
    outputs(6818) <= not(layer2_outputs(4687));
    outputs(6819) <= layer2_outputs(8884);
    outputs(6820) <= not((layer2_outputs(8437)) xor (layer2_outputs(2993)));
    outputs(6821) <= not(layer2_outputs(361));
    outputs(6822) <= not(layer2_outputs(2444));
    outputs(6823) <= not(layer2_outputs(7341));
    outputs(6824) <= not(layer2_outputs(2033));
    outputs(6825) <= (layer2_outputs(1931)) xor (layer2_outputs(5260));
    outputs(6826) <= not(layer2_outputs(4009));
    outputs(6827) <= layer2_outputs(7692);
    outputs(6828) <= not(layer2_outputs(7083));
    outputs(6829) <= layer2_outputs(2439);
    outputs(6830) <= not(layer2_outputs(4807));
    outputs(6831) <= not(layer2_outputs(8073));
    outputs(6832) <= not(layer2_outputs(252));
    outputs(6833) <= not(layer2_outputs(4839));
    outputs(6834) <= layer2_outputs(7455);
    outputs(6835) <= not(layer2_outputs(2791));
    outputs(6836) <= layer2_outputs(7768);
    outputs(6837) <= not(layer2_outputs(240));
    outputs(6838) <= not(layer2_outputs(5054));
    outputs(6839) <= not((layer2_outputs(6085)) xor (layer2_outputs(4545)));
    outputs(6840) <= layer2_outputs(1338);
    outputs(6841) <= not(layer2_outputs(1504));
    outputs(6842) <= layer2_outputs(2135);
    outputs(6843) <= (layer2_outputs(272)) and not (layer2_outputs(7224));
    outputs(6844) <= layer2_outputs(9477);
    outputs(6845) <= (layer2_outputs(126)) and not (layer2_outputs(6846));
    outputs(6846) <= (layer2_outputs(2615)) and not (layer2_outputs(3245));
    outputs(6847) <= not(layer2_outputs(9099));
    outputs(6848) <= not((layer2_outputs(1091)) xor (layer2_outputs(8518)));
    outputs(6849) <= layer2_outputs(4004);
    outputs(6850) <= not(layer2_outputs(4561));
    outputs(6851) <= (layer2_outputs(501)) and not (layer2_outputs(398));
    outputs(6852) <= not(layer2_outputs(2027));
    outputs(6853) <= layer2_outputs(7639);
    outputs(6854) <= not(layer2_outputs(2809));
    outputs(6855) <= not((layer2_outputs(3431)) xor (layer2_outputs(3224)));
    outputs(6856) <= not((layer2_outputs(8950)) xor (layer2_outputs(954)));
    outputs(6857) <= not((layer2_outputs(10211)) or (layer2_outputs(6983)));
    outputs(6858) <= (layer2_outputs(64)) and not (layer2_outputs(9760));
    outputs(6859) <= (layer2_outputs(983)) xor (layer2_outputs(2022));
    outputs(6860) <= (layer2_outputs(6534)) xor (layer2_outputs(4780));
    outputs(6861) <= (layer2_outputs(5174)) xor (layer2_outputs(5343));
    outputs(6862) <= not((layer2_outputs(371)) xor (layer2_outputs(7948)));
    outputs(6863) <= not(layer2_outputs(5584));
    outputs(6864) <= not(layer2_outputs(7557));
    outputs(6865) <= layer2_outputs(7769);
    outputs(6866) <= not(layer2_outputs(8149));
    outputs(6867) <= (layer2_outputs(8638)) and (layer2_outputs(2199));
    outputs(6868) <= layer2_outputs(2510);
    outputs(6869) <= layer2_outputs(8834);
    outputs(6870) <= not(layer2_outputs(7289));
    outputs(6871) <= not(layer2_outputs(4835)) or (layer2_outputs(6144));
    outputs(6872) <= layer2_outputs(3259);
    outputs(6873) <= layer2_outputs(2555);
    outputs(6874) <= not(layer2_outputs(1313));
    outputs(6875) <= not(layer2_outputs(2862));
    outputs(6876) <= (layer2_outputs(7869)) xor (layer2_outputs(1784));
    outputs(6877) <= not(layer2_outputs(6975));
    outputs(6878) <= not((layer2_outputs(1085)) or (layer2_outputs(3659)));
    outputs(6879) <= not((layer2_outputs(9372)) or (layer2_outputs(6160)));
    outputs(6880) <= not(layer2_outputs(9479));
    outputs(6881) <= not(layer2_outputs(3793));
    outputs(6882) <= not((layer2_outputs(5547)) or (layer2_outputs(7698)));
    outputs(6883) <= not(layer2_outputs(9310));
    outputs(6884) <= layer2_outputs(6406);
    outputs(6885) <= not((layer2_outputs(8676)) and (layer2_outputs(2768)));
    outputs(6886) <= not(layer2_outputs(3619));
    outputs(6887) <= not((layer2_outputs(3406)) xor (layer2_outputs(5243)));
    outputs(6888) <= not(layer2_outputs(4239));
    outputs(6889) <= not((layer2_outputs(8186)) or (layer2_outputs(9211)));
    outputs(6890) <= layer2_outputs(7604);
    outputs(6891) <= layer2_outputs(1794);
    outputs(6892) <= not(layer2_outputs(5701));
    outputs(6893) <= layer2_outputs(2331);
    outputs(6894) <= layer2_outputs(7352);
    outputs(6895) <= layer2_outputs(9741);
    outputs(6896) <= not(layer2_outputs(3668));
    outputs(6897) <= not(layer2_outputs(7269));
    outputs(6898) <= not((layer2_outputs(6752)) xor (layer2_outputs(5029)));
    outputs(6899) <= not(layer2_outputs(1276));
    outputs(6900) <= not(layer2_outputs(1705));
    outputs(6901) <= (layer2_outputs(1901)) xor (layer2_outputs(7362));
    outputs(6902) <= not(layer2_outputs(2163));
    outputs(6903) <= not(layer2_outputs(9385));
    outputs(6904) <= (layer2_outputs(3456)) and not (layer2_outputs(9120));
    outputs(6905) <= not(layer2_outputs(9377));
    outputs(6906) <= layer2_outputs(7974);
    outputs(6907) <= not(layer2_outputs(2740)) or (layer2_outputs(9386));
    outputs(6908) <= not(layer2_outputs(9886));
    outputs(6909) <= layer2_outputs(1801);
    outputs(6910) <= layer2_outputs(5906);
    outputs(6911) <= not((layer2_outputs(3055)) xor (layer2_outputs(9614)));
    outputs(6912) <= layer2_outputs(3968);
    outputs(6913) <= layer2_outputs(7003);
    outputs(6914) <= not(layer2_outputs(5429));
    outputs(6915) <= layer2_outputs(3876);
    outputs(6916) <= (layer2_outputs(4785)) xor (layer2_outputs(6121));
    outputs(6917) <= not(layer2_outputs(6085));
    outputs(6918) <= layer2_outputs(8700);
    outputs(6919) <= layer2_outputs(1879);
    outputs(6920) <= (layer2_outputs(8908)) xor (layer2_outputs(10025));
    outputs(6921) <= (layer2_outputs(7331)) and not (layer2_outputs(7089));
    outputs(6922) <= not(layer2_outputs(4839)) or (layer2_outputs(6512));
    outputs(6923) <= (layer2_outputs(2544)) xor (layer2_outputs(4947));
    outputs(6924) <= layer2_outputs(9264);
    outputs(6925) <= layer2_outputs(3069);
    outputs(6926) <= not(layer2_outputs(8522));
    outputs(6927) <= layer2_outputs(2595);
    outputs(6928) <= not(layer2_outputs(4883));
    outputs(6929) <= layer2_outputs(2755);
    outputs(6930) <= not(layer2_outputs(9318));
    outputs(6931) <= layer2_outputs(8759);
    outputs(6932) <= not((layer2_outputs(9649)) xor (layer2_outputs(4206)));
    outputs(6933) <= layer2_outputs(6363);
    outputs(6934) <= not(layer2_outputs(5675));
    outputs(6935) <= not(layer2_outputs(6194));
    outputs(6936) <= not((layer2_outputs(1279)) or (layer2_outputs(9625)));
    outputs(6937) <= layer2_outputs(6167);
    outputs(6938) <= not(layer2_outputs(3510));
    outputs(6939) <= not(layer2_outputs(6225));
    outputs(6940) <= not(layer2_outputs(9574));
    outputs(6941) <= layer2_outputs(2792);
    outputs(6942) <= layer2_outputs(388);
    outputs(6943) <= layer2_outputs(6465);
    outputs(6944) <= layer2_outputs(5111);
    outputs(6945) <= not(layer2_outputs(2789));
    outputs(6946) <= layer2_outputs(5567);
    outputs(6947) <= not(layer2_outputs(8137)) or (layer2_outputs(4179));
    outputs(6948) <= layer2_outputs(7380);
    outputs(6949) <= not(layer2_outputs(7457));
    outputs(6950) <= layer2_outputs(5182);
    outputs(6951) <= not(layer2_outputs(5297));
    outputs(6952) <= not(layer2_outputs(8996));
    outputs(6953) <= not(layer2_outputs(976));
    outputs(6954) <= not((layer2_outputs(6521)) xor (layer2_outputs(8764)));
    outputs(6955) <= layer2_outputs(2833);
    outputs(6956) <= (layer2_outputs(1244)) and not (layer2_outputs(3286));
    outputs(6957) <= not(layer2_outputs(8012));
    outputs(6958) <= not(layer2_outputs(4252));
    outputs(6959) <= not(layer2_outputs(3228));
    outputs(6960) <= layer2_outputs(8128);
    outputs(6961) <= not(layer2_outputs(1482));
    outputs(6962) <= not((layer2_outputs(160)) xor (layer2_outputs(6270)));
    outputs(6963) <= layer2_outputs(7248);
    outputs(6964) <= layer2_outputs(4109);
    outputs(6965) <= not(layer2_outputs(1656));
    outputs(6966) <= (layer2_outputs(7432)) xor (layer2_outputs(6336));
    outputs(6967) <= layer2_outputs(3016);
    outputs(6968) <= layer2_outputs(3603);
    outputs(6969) <= not(layer2_outputs(9357));
    outputs(6970) <= layer2_outputs(7497);
    outputs(6971) <= (layer2_outputs(50)) and not (layer2_outputs(8075));
    outputs(6972) <= layer2_outputs(9198);
    outputs(6973) <= layer2_outputs(5568);
    outputs(6974) <= layer2_outputs(6044);
    outputs(6975) <= layer2_outputs(7801);
    outputs(6976) <= layer2_outputs(2554);
    outputs(6977) <= (layer2_outputs(4000)) and not (layer2_outputs(7190));
    outputs(6978) <= not(layer2_outputs(7421));
    outputs(6979) <= not(layer2_outputs(6128));
    outputs(6980) <= layer2_outputs(253);
    outputs(6981) <= layer2_outputs(675);
    outputs(6982) <= not((layer2_outputs(9101)) or (layer2_outputs(6104)));
    outputs(6983) <= layer2_outputs(10064);
    outputs(6984) <= layer2_outputs(3069);
    outputs(6985) <= (layer2_outputs(8124)) and (layer2_outputs(1941));
    outputs(6986) <= layer2_outputs(8414);
    outputs(6987) <= not((layer2_outputs(3096)) xor (layer2_outputs(3854)));
    outputs(6988) <= not(layer2_outputs(7084));
    outputs(6989) <= not(layer2_outputs(7124));
    outputs(6990) <= not(layer2_outputs(3250));
    outputs(6991) <= not(layer2_outputs(706));
    outputs(6992) <= (layer2_outputs(7773)) xor (layer2_outputs(3024));
    outputs(6993) <= (layer2_outputs(4856)) xor (layer2_outputs(5507));
    outputs(6994) <= layer2_outputs(5740);
    outputs(6995) <= not(layer2_outputs(2668));
    outputs(6996) <= not((layer2_outputs(4938)) xor (layer2_outputs(6631)));
    outputs(6997) <= layer2_outputs(9459);
    outputs(6998) <= not(layer2_outputs(2136));
    outputs(6999) <= (layer2_outputs(8216)) and not (layer2_outputs(5430));
    outputs(7000) <= layer2_outputs(10141);
    outputs(7001) <= not((layer2_outputs(4170)) xor (layer2_outputs(179)));
    outputs(7002) <= layer2_outputs(3203);
    outputs(7003) <= layer2_outputs(5225);
    outputs(7004) <= layer2_outputs(9642);
    outputs(7005) <= not(layer2_outputs(251)) or (layer2_outputs(10168));
    outputs(7006) <= layer2_outputs(1440);
    outputs(7007) <= layer2_outputs(5930);
    outputs(7008) <= layer2_outputs(8138);
    outputs(7009) <= layer2_outputs(8144);
    outputs(7010) <= (layer2_outputs(7791)) and (layer2_outputs(44));
    outputs(7011) <= (layer2_outputs(7940)) and not (layer2_outputs(7491));
    outputs(7012) <= not(layer2_outputs(6082));
    outputs(7013) <= layer2_outputs(3615);
    outputs(7014) <= layer2_outputs(8345);
    outputs(7015) <= not(layer2_outputs(8451));
    outputs(7016) <= (layer2_outputs(6032)) and not (layer2_outputs(1923));
    outputs(7017) <= layer2_outputs(760);
    outputs(7018) <= layer2_outputs(3803);
    outputs(7019) <= (layer2_outputs(6853)) xor (layer2_outputs(4677));
    outputs(7020) <= layer2_outputs(8401);
    outputs(7021) <= layer2_outputs(591);
    outputs(7022) <= layer2_outputs(5549);
    outputs(7023) <= (layer2_outputs(3441)) xor (layer2_outputs(832));
    outputs(7024) <= (layer2_outputs(1664)) and (layer2_outputs(2165));
    outputs(7025) <= layer2_outputs(3781);
    outputs(7026) <= not((layer2_outputs(2089)) xor (layer2_outputs(3289)));
    outputs(7027) <= not((layer2_outputs(6499)) xor (layer2_outputs(6938)));
    outputs(7028) <= not(layer2_outputs(3127));
    outputs(7029) <= layer2_outputs(4531);
    outputs(7030) <= layer2_outputs(4158);
    outputs(7031) <= not(layer2_outputs(1212));
    outputs(7032) <= layer2_outputs(6756);
    outputs(7033) <= layer2_outputs(2542);
    outputs(7034) <= (layer2_outputs(6031)) xor (layer2_outputs(6826));
    outputs(7035) <= not((layer2_outputs(7594)) xor (layer2_outputs(8341)));
    outputs(7036) <= layer2_outputs(5549);
    outputs(7037) <= layer2_outputs(7598);
    outputs(7038) <= layer2_outputs(1939);
    outputs(7039) <= (layer2_outputs(9907)) and (layer2_outputs(1419));
    outputs(7040) <= layer2_outputs(3442);
    outputs(7041) <= layer2_outputs(563);
    outputs(7042) <= (layer2_outputs(1035)) xor (layer2_outputs(8146));
    outputs(7043) <= layer2_outputs(1385);
    outputs(7044) <= not(layer2_outputs(9927));
    outputs(7045) <= (layer2_outputs(7691)) and (layer2_outputs(3828));
    outputs(7046) <= not((layer2_outputs(4559)) xor (layer2_outputs(1042)));
    outputs(7047) <= not(layer2_outputs(1019));
    outputs(7048) <= (layer2_outputs(3874)) xor (layer2_outputs(1917));
    outputs(7049) <= layer2_outputs(10149);
    outputs(7050) <= not(layer2_outputs(6808));
    outputs(7051) <= not((layer2_outputs(8521)) or (layer2_outputs(3122)));
    outputs(7052) <= not((layer2_outputs(4308)) and (layer2_outputs(4463)));
    outputs(7053) <= not((layer2_outputs(6735)) or (layer2_outputs(3108)));
    outputs(7054) <= (layer2_outputs(9602)) xor (layer2_outputs(3787));
    outputs(7055) <= not((layer2_outputs(9807)) and (layer2_outputs(4781)));
    outputs(7056) <= not((layer2_outputs(3535)) xor (layer2_outputs(2264)));
    outputs(7057) <= layer2_outputs(7809);
    outputs(7058) <= (layer2_outputs(6294)) xor (layer2_outputs(5552));
    outputs(7059) <= (layer2_outputs(9710)) and not (layer2_outputs(6023));
    outputs(7060) <= layer2_outputs(5313);
    outputs(7061) <= layer2_outputs(8360);
    outputs(7062) <= not(layer2_outputs(6661));
    outputs(7063) <= (layer2_outputs(6493)) xor (layer2_outputs(6238));
    outputs(7064) <= not((layer2_outputs(5639)) and (layer2_outputs(2929)));
    outputs(7065) <= layer2_outputs(8514);
    outputs(7066) <= layer2_outputs(6289);
    outputs(7067) <= (layer2_outputs(7898)) xor (layer2_outputs(9506));
    outputs(7068) <= layer2_outputs(2856);
    outputs(7069) <= not(layer2_outputs(1753));
    outputs(7070) <= (layer2_outputs(1426)) and not (layer2_outputs(5943));
    outputs(7071) <= not(layer2_outputs(4393));
    outputs(7072) <= layer2_outputs(3022);
    outputs(7073) <= not(layer2_outputs(1175));
    outputs(7074) <= not((layer2_outputs(5369)) or (layer2_outputs(7062)));
    outputs(7075) <= layer2_outputs(3561);
    outputs(7076) <= not(layer2_outputs(262));
    outputs(7077) <= (layer2_outputs(222)) and not (layer2_outputs(1678));
    outputs(7078) <= not(layer2_outputs(1911));
    outputs(7079) <= (layer2_outputs(2056)) and not (layer2_outputs(5181));
    outputs(7080) <= layer2_outputs(5171);
    outputs(7081) <= layer2_outputs(9984);
    outputs(7082) <= not(layer2_outputs(217));
    outputs(7083) <= not(layer2_outputs(789));
    outputs(7084) <= not(layer2_outputs(8166)) or (layer2_outputs(3866));
    outputs(7085) <= not(layer2_outputs(9820));
    outputs(7086) <= layer2_outputs(3518);
    outputs(7087) <= not((layer2_outputs(2018)) xor (layer2_outputs(4975)));
    outputs(7088) <= not((layer2_outputs(6613)) and (layer2_outputs(5954)));
    outputs(7089) <= (layer2_outputs(6468)) and not (layer2_outputs(4991));
    outputs(7090) <= layer2_outputs(9187);
    outputs(7091) <= layer2_outputs(8848);
    outputs(7092) <= (layer2_outputs(2328)) xor (layer2_outputs(2956));
    outputs(7093) <= (layer2_outputs(3056)) or (layer2_outputs(6711));
    outputs(7094) <= layer2_outputs(8800);
    outputs(7095) <= (layer2_outputs(4062)) and (layer2_outputs(9171));
    outputs(7096) <= not(layer2_outputs(4568));
    outputs(7097) <= not(layer2_outputs(6060));
    outputs(7098) <= layer2_outputs(10048);
    outputs(7099) <= not(layer2_outputs(165));
    outputs(7100) <= layer2_outputs(5940);
    outputs(7101) <= layer2_outputs(1099);
    outputs(7102) <= layer2_outputs(3386);
    outputs(7103) <= not(layer2_outputs(366));
    outputs(7104) <= not(layer2_outputs(4210));
    outputs(7105) <= (layer2_outputs(4060)) and (layer2_outputs(4191));
    outputs(7106) <= (layer2_outputs(8630)) xor (layer2_outputs(756));
    outputs(7107) <= not(layer2_outputs(1841));
    outputs(7108) <= not(layer2_outputs(8467));
    outputs(7109) <= layer2_outputs(4294);
    outputs(7110) <= (layer2_outputs(1012)) and not (layer2_outputs(6871));
    outputs(7111) <= (layer2_outputs(2816)) xor (layer2_outputs(7985));
    outputs(7112) <= not(layer2_outputs(9812));
    outputs(7113) <= layer2_outputs(10124);
    outputs(7114) <= not((layer2_outputs(9224)) or (layer2_outputs(1038)));
    outputs(7115) <= not(layer2_outputs(9482));
    outputs(7116) <= (layer2_outputs(8308)) and not (layer2_outputs(242));
    outputs(7117) <= not((layer2_outputs(2371)) xor (layer2_outputs(7584)));
    outputs(7118) <= (layer2_outputs(8868)) xor (layer2_outputs(2646));
    outputs(7119) <= not(layer2_outputs(5869)) or (layer2_outputs(2074));
    outputs(7120) <= layer2_outputs(781);
    outputs(7121) <= not((layer2_outputs(9536)) xor (layer2_outputs(8416)));
    outputs(7122) <= layer2_outputs(2636);
    outputs(7123) <= not(layer2_outputs(9923));
    outputs(7124) <= not(layer2_outputs(9382));
    outputs(7125) <= not(layer2_outputs(9750)) or (layer2_outputs(3193));
    outputs(7126) <= not(layer2_outputs(3830));
    outputs(7127) <= layer2_outputs(1922);
    outputs(7128) <= not((layer2_outputs(3964)) xor (layer2_outputs(72)));
    outputs(7129) <= not((layer2_outputs(6234)) xor (layer2_outputs(9861)));
    outputs(7130) <= (layer2_outputs(2469)) xor (layer2_outputs(4706));
    outputs(7131) <= not((layer2_outputs(5478)) xor (layer2_outputs(6344)));
    outputs(7132) <= not((layer2_outputs(208)) or (layer2_outputs(8844)));
    outputs(7133) <= not(layer2_outputs(554));
    outputs(7134) <= layer2_outputs(3533);
    outputs(7135) <= not(layer2_outputs(3144));
    outputs(7136) <= layer2_outputs(9337);
    outputs(7137) <= (layer2_outputs(6705)) and not (layer2_outputs(6848));
    outputs(7138) <= not(layer2_outputs(9144));
    outputs(7139) <= (layer2_outputs(2595)) and not (layer2_outputs(8656));
    outputs(7140) <= (layer2_outputs(1566)) or (layer2_outputs(8991));
    outputs(7141) <= (layer2_outputs(3750)) xor (layer2_outputs(5638));
    outputs(7142) <= not(layer2_outputs(2132));
    outputs(7143) <= not(layer2_outputs(5994));
    outputs(7144) <= not((layer2_outputs(1161)) xor (layer2_outputs(9030)));
    outputs(7145) <= not(layer2_outputs(3312));
    outputs(7146) <= layer2_outputs(2142);
    outputs(7147) <= not(layer2_outputs(5717));
    outputs(7148) <= not(layer2_outputs(5304)) or (layer2_outputs(8389));
    outputs(7149) <= layer2_outputs(4342);
    outputs(7150) <= not(layer2_outputs(5929)) or (layer2_outputs(1320));
    outputs(7151) <= (layer2_outputs(7967)) xor (layer2_outputs(1289));
    outputs(7152) <= layer2_outputs(2629);
    outputs(7153) <= not(layer2_outputs(5898));
    outputs(7154) <= not(layer2_outputs(4301));
    outputs(7155) <= layer2_outputs(8498);
    outputs(7156) <= layer2_outputs(351);
    outputs(7157) <= not(layer2_outputs(2303));
    outputs(7158) <= not(layer2_outputs(5361));
    outputs(7159) <= layer2_outputs(5723);
    outputs(7160) <= layer2_outputs(8943);
    outputs(7161) <= (layer2_outputs(1134)) and not (layer2_outputs(1691));
    outputs(7162) <= layer2_outputs(3782);
    outputs(7163) <= layer2_outputs(9304);
    outputs(7164) <= layer2_outputs(7516);
    outputs(7165) <= layer2_outputs(1496);
    outputs(7166) <= layer2_outputs(1900);
    outputs(7167) <= layer2_outputs(4637);
    outputs(7168) <= (layer2_outputs(3982)) and not (layer2_outputs(1292));
    outputs(7169) <= layer2_outputs(4821);
    outputs(7170) <= not(layer2_outputs(3577));
    outputs(7171) <= layer2_outputs(8556);
    outputs(7172) <= layer2_outputs(5275);
    outputs(7173) <= not(layer2_outputs(7747));
    outputs(7174) <= not(layer2_outputs(148));
    outputs(7175) <= not(layer2_outputs(4045));
    outputs(7176) <= layer2_outputs(4533);
    outputs(7177) <= not(layer2_outputs(2190)) or (layer2_outputs(1523));
    outputs(7178) <= not(layer2_outputs(9443));
    outputs(7179) <= not(layer2_outputs(4127));
    outputs(7180) <= layer2_outputs(1497);
    outputs(7181) <= not(layer2_outputs(5290));
    outputs(7182) <= (layer2_outputs(6608)) and not (layer2_outputs(9151));
    outputs(7183) <= not((layer2_outputs(3802)) xor (layer2_outputs(1438)));
    outputs(7184) <= layer2_outputs(4068);
    outputs(7185) <= layer2_outputs(7290);
    outputs(7186) <= (layer2_outputs(1948)) and not (layer2_outputs(3076));
    outputs(7187) <= (layer2_outputs(224)) or (layer2_outputs(2456));
    outputs(7188) <= not(layer2_outputs(5661));
    outputs(7189) <= layer2_outputs(2657);
    outputs(7190) <= layer2_outputs(926);
    outputs(7191) <= not(layer2_outputs(8480));
    outputs(7192) <= not(layer2_outputs(9631));
    outputs(7193) <= (layer2_outputs(580)) xor (layer2_outputs(8220));
    outputs(7194) <= not((layer2_outputs(4629)) or (layer2_outputs(3081)));
    outputs(7195) <= not((layer2_outputs(3817)) xor (layer2_outputs(3564)));
    outputs(7196) <= (layer2_outputs(1568)) and not (layer2_outputs(1219));
    outputs(7197) <= (layer2_outputs(5115)) xor (layer2_outputs(2827));
    outputs(7198) <= layer2_outputs(6528);
    outputs(7199) <= layer2_outputs(8934);
    outputs(7200) <= not(layer2_outputs(4173));
    outputs(7201) <= not((layer2_outputs(7474)) or (layer2_outputs(561)));
    outputs(7202) <= not(layer2_outputs(1903));
    outputs(7203) <= not(layer2_outputs(10185));
    outputs(7204) <= layer2_outputs(5767);
    outputs(7205) <= not((layer2_outputs(3045)) xor (layer2_outputs(2338)));
    outputs(7206) <= not((layer2_outputs(1475)) xor (layer2_outputs(1919)));
    outputs(7207) <= (layer2_outputs(6147)) xor (layer2_outputs(9271));
    outputs(7208) <= (layer2_outputs(3350)) and not (layer2_outputs(661));
    outputs(7209) <= not(layer2_outputs(8512));
    outputs(7210) <= layer2_outputs(9483);
    outputs(7211) <= not(layer2_outputs(7129)) or (layer2_outputs(1977));
    outputs(7212) <= not(layer2_outputs(6543));
    outputs(7213) <= layer2_outputs(7290);
    outputs(7214) <= layer2_outputs(845);
    outputs(7215) <= not(layer2_outputs(1189)) or (layer2_outputs(10146));
    outputs(7216) <= not((layer2_outputs(8767)) or (layer2_outputs(8364)));
    outputs(7217) <= layer2_outputs(1815);
    outputs(7218) <= layer2_outputs(1655);
    outputs(7219) <= layer2_outputs(4418);
    outputs(7220) <= layer2_outputs(5539);
    outputs(7221) <= not(layer2_outputs(1754));
    outputs(7222) <= layer2_outputs(2303);
    outputs(7223) <= not(layer2_outputs(3590));
    outputs(7224) <= not(layer2_outputs(3193));
    outputs(7225) <= (layer2_outputs(8245)) and not (layer2_outputs(1659));
    outputs(7226) <= layer2_outputs(7895);
    outputs(7227) <= layer2_outputs(3959);
    outputs(7228) <= not(layer2_outputs(8344));
    outputs(7229) <= not(layer2_outputs(1515));
    outputs(7230) <= layer2_outputs(9024);
    outputs(7231) <= layer2_outputs(559);
    outputs(7232) <= not((layer2_outputs(10155)) xor (layer2_outputs(9266)));
    outputs(7233) <= not(layer2_outputs(5428));
    outputs(7234) <= (layer2_outputs(9012)) and not (layer2_outputs(4689));
    outputs(7235) <= not(layer2_outputs(2200));
    outputs(7236) <= not(layer2_outputs(3229));
    outputs(7237) <= not(layer2_outputs(8143)) or (layer2_outputs(885));
    outputs(7238) <= not(layer2_outputs(6092));
    outputs(7239) <= not(layer2_outputs(112));
    outputs(7240) <= layer2_outputs(2617);
    outputs(7241) <= layer2_outputs(8963);
    outputs(7242) <= (layer2_outputs(5461)) xor (layer2_outputs(8488));
    outputs(7243) <= (layer2_outputs(6196)) and not (layer2_outputs(7093));
    outputs(7244) <= not(layer2_outputs(4384));
    outputs(7245) <= not(layer2_outputs(921));
    outputs(7246) <= layer2_outputs(327);
    outputs(7247) <= layer2_outputs(2092);
    outputs(7248) <= (layer2_outputs(7414)) and not (layer2_outputs(9118));
    outputs(7249) <= not((layer2_outputs(4611)) or (layer2_outputs(2124)));
    outputs(7250) <= not(layer2_outputs(4151));
    outputs(7251) <= layer2_outputs(5305);
    outputs(7252) <= layer2_outputs(3134);
    outputs(7253) <= layer2_outputs(1891);
    outputs(7254) <= layer2_outputs(7089);
    outputs(7255) <= (layer2_outputs(8533)) xor (layer2_outputs(570));
    outputs(7256) <= not(layer2_outputs(7208)) or (layer2_outputs(1534));
    outputs(7257) <= layer2_outputs(9201);
    outputs(7258) <= not(layer2_outputs(2278));
    outputs(7259) <= layer2_outputs(8166);
    outputs(7260) <= (layer2_outputs(9312)) xor (layer2_outputs(6337));
    outputs(7261) <= not(layer2_outputs(1547));
    outputs(7262) <= layer2_outputs(6243);
    outputs(7263) <= layer2_outputs(1116);
    outputs(7264) <= layer2_outputs(7568);
    outputs(7265) <= not((layer2_outputs(917)) or (layer2_outputs(1430)));
    outputs(7266) <= not(layer2_outputs(8608));
    outputs(7267) <= (layer2_outputs(1444)) xor (layer2_outputs(1915));
    outputs(7268) <= not(layer2_outputs(7581));
    outputs(7269) <= layer2_outputs(4925);
    outputs(7270) <= not((layer2_outputs(4920)) and (layer2_outputs(5086)));
    outputs(7271) <= layer2_outputs(1815);
    outputs(7272) <= not(layer2_outputs(6069));
    outputs(7273) <= not(layer2_outputs(1851));
    outputs(7274) <= (layer2_outputs(5726)) and (layer2_outputs(7741));
    outputs(7275) <= layer2_outputs(2414);
    outputs(7276) <= not(layer2_outputs(4093));
    outputs(7277) <= layer2_outputs(7049);
    outputs(7278) <= (layer2_outputs(313)) xor (layer2_outputs(1150));
    outputs(7279) <= not(layer2_outputs(8040));
    outputs(7280) <= layer2_outputs(9132);
    outputs(7281) <= layer2_outputs(671);
    outputs(7282) <= (layer2_outputs(3550)) and not (layer2_outputs(9896));
    outputs(7283) <= not(layer2_outputs(7077));
    outputs(7284) <= not(layer2_outputs(7323));
    outputs(7285) <= not(layer2_outputs(7199)) or (layer2_outputs(3679));
    outputs(7286) <= (layer2_outputs(6202)) and not (layer2_outputs(8670));
    outputs(7287) <= layer2_outputs(859);
    outputs(7288) <= layer2_outputs(5450);
    outputs(7289) <= not((layer2_outputs(7326)) xor (layer2_outputs(2532)));
    outputs(7290) <= not(layer2_outputs(6561));
    outputs(7291) <= (layer2_outputs(522)) and not (layer2_outputs(4956));
    outputs(7292) <= (layer2_outputs(9123)) and (layer2_outputs(2041));
    outputs(7293) <= not(layer2_outputs(2116));
    outputs(7294) <= not(layer2_outputs(1747));
    outputs(7295) <= (layer2_outputs(3358)) and (layer2_outputs(1003));
    outputs(7296) <= not(layer2_outputs(8279));
    outputs(7297) <= not((layer2_outputs(9944)) or (layer2_outputs(3798)));
    outputs(7298) <= not(layer2_outputs(8485));
    outputs(7299) <= layer2_outputs(4128);
    outputs(7300) <= (layer2_outputs(2292)) xor (layer2_outputs(5380));
    outputs(7301) <= layer2_outputs(7127);
    outputs(7302) <= layer2_outputs(8579);
    outputs(7303) <= not(layer2_outputs(6833));
    outputs(7304) <= layer2_outputs(4575);
    outputs(7305) <= layer2_outputs(1178);
    outputs(7306) <= (layer2_outputs(3377)) and not (layer2_outputs(828));
    outputs(7307) <= not((layer2_outputs(3394)) xor (layer2_outputs(8125)));
    outputs(7308) <= not((layer2_outputs(4918)) xor (layer2_outputs(7331)));
    outputs(7309) <= not(layer2_outputs(3970));
    outputs(7310) <= (layer2_outputs(5089)) xor (layer2_outputs(7605));
    outputs(7311) <= layer2_outputs(774);
    outputs(7312) <= (layer2_outputs(947)) and not (layer2_outputs(6847));
    outputs(7313) <= (layer2_outputs(5916)) and (layer2_outputs(6649));
    outputs(7314) <= not(layer2_outputs(9461));
    outputs(7315) <= layer2_outputs(7471);
    outputs(7316) <= not(layer2_outputs(6766));
    outputs(7317) <= not(layer2_outputs(761)) or (layer2_outputs(7520));
    outputs(7318) <= (layer2_outputs(5222)) and (layer2_outputs(5869));
    outputs(7319) <= layer2_outputs(9338);
    outputs(7320) <= (layer2_outputs(1899)) xor (layer2_outputs(736));
    outputs(7321) <= layer2_outputs(3083);
    outputs(7322) <= layer2_outputs(2650);
    outputs(7323) <= not((layer2_outputs(10120)) or (layer2_outputs(6405)));
    outputs(7324) <= (layer2_outputs(5530)) and not (layer2_outputs(5859));
    outputs(7325) <= not(layer2_outputs(3313));
    outputs(7326) <= (layer2_outputs(6036)) xor (layer2_outputs(3829));
    outputs(7327) <= not((layer2_outputs(6058)) xor (layer2_outputs(6115)));
    outputs(7328) <= (layer2_outputs(8464)) and (layer2_outputs(10017));
    outputs(7329) <= not(layer2_outputs(5999));
    outputs(7330) <= layer2_outputs(1834);
    outputs(7331) <= layer2_outputs(7492);
    outputs(7332) <= not(layer2_outputs(4886));
    outputs(7333) <= not(layer2_outputs(5357));
    outputs(7334) <= not((layer2_outputs(4751)) xor (layer2_outputs(5603)));
    outputs(7335) <= not(layer2_outputs(4114));
    outputs(7336) <= layer2_outputs(8173);
    outputs(7337) <= layer2_outputs(1686);
    outputs(7338) <= layer2_outputs(4415);
    outputs(7339) <= not(layer2_outputs(299));
    outputs(7340) <= not(layer2_outputs(669));
    outputs(7341) <= layer2_outputs(6302);
    outputs(7342) <= not(layer2_outputs(1002));
    outputs(7343) <= not((layer2_outputs(8785)) and (layer2_outputs(5565)));
    outputs(7344) <= (layer2_outputs(10037)) and not (layer2_outputs(3566));
    outputs(7345) <= layer2_outputs(8121);
    outputs(7346) <= layer2_outputs(10050);
    outputs(7347) <= (layer2_outputs(4374)) xor (layer2_outputs(7535));
    outputs(7348) <= (layer2_outputs(1512)) or (layer2_outputs(8187));
    outputs(7349) <= not(layer2_outputs(6215));
    outputs(7350) <= not(layer2_outputs(2076)) or (layer2_outputs(3625));
    outputs(7351) <= not((layer2_outputs(126)) or (layer2_outputs(9167)));
    outputs(7352) <= not((layer2_outputs(1201)) xor (layer2_outputs(1570)));
    outputs(7353) <= (layer2_outputs(8202)) and (layer2_outputs(3674));
    outputs(7354) <= not(layer2_outputs(8155));
    outputs(7355) <= (layer2_outputs(246)) and not (layer2_outputs(5968));
    outputs(7356) <= not(layer2_outputs(649));
    outputs(7357) <= not(layer2_outputs(6676));
    outputs(7358) <= layer2_outputs(448);
    outputs(7359) <= (layer2_outputs(5805)) and (layer2_outputs(3408));
    outputs(7360) <= layer2_outputs(4232);
    outputs(7361) <= layer2_outputs(3465);
    outputs(7362) <= not(layer2_outputs(962));
    outputs(7363) <= layer2_outputs(7602);
    outputs(7364) <= not(layer2_outputs(6407));
    outputs(7365) <= not(layer2_outputs(6321));
    outputs(7366) <= layer2_outputs(5301);
    outputs(7367) <= not(layer2_outputs(6764));
    outputs(7368) <= (layer2_outputs(1994)) xor (layer2_outputs(2725));
    outputs(7369) <= layer2_outputs(5402);
    outputs(7370) <= layer2_outputs(721);
    outputs(7371) <= layer2_outputs(4460);
    outputs(7372) <= layer2_outputs(7448);
    outputs(7373) <= not(layer2_outputs(4215));
    outputs(7374) <= layer2_outputs(7101);
    outputs(7375) <= not(layer2_outputs(7305));
    outputs(7376) <= (layer2_outputs(9806)) xor (layer2_outputs(3017));
    outputs(7377) <= layer2_outputs(6945);
    outputs(7378) <= not(layer2_outputs(8902));
    outputs(7379) <= not((layer2_outputs(982)) xor (layer2_outputs(7432)));
    outputs(7380) <= layer2_outputs(2046);
    outputs(7381) <= layer2_outputs(3523);
    outputs(7382) <= not(layer2_outputs(6770));
    outputs(7383) <= not(layer2_outputs(1680));
    outputs(7384) <= not(layer2_outputs(8127));
    outputs(7385) <= (layer2_outputs(4482)) xor (layer2_outputs(8037));
    outputs(7386) <= not((layer2_outputs(4141)) xor (layer2_outputs(8333)));
    outputs(7387) <= not((layer2_outputs(9199)) or (layer2_outputs(5320)));
    outputs(7388) <= layer2_outputs(8171);
    outputs(7389) <= not((layer2_outputs(7094)) xor (layer2_outputs(5564)));
    outputs(7390) <= layer2_outputs(6699);
    outputs(7391) <= not(layer2_outputs(8563));
    outputs(7392) <= not(layer2_outputs(3822));
    outputs(7393) <= layer2_outputs(4242);
    outputs(7394) <= (layer2_outputs(4757)) and not (layer2_outputs(6559));
    outputs(7395) <= not(layer2_outputs(3764));
    outputs(7396) <= layer2_outputs(6828);
    outputs(7397) <= (layer2_outputs(8103)) and not (layer2_outputs(7783));
    outputs(7398) <= (layer2_outputs(6008)) xor (layer2_outputs(2665));
    outputs(7399) <= layer2_outputs(4029);
    outputs(7400) <= not(layer2_outputs(2315));
    outputs(7401) <= (layer2_outputs(10207)) and not (layer2_outputs(6236));
    outputs(7402) <= layer2_outputs(2539);
    outputs(7403) <= layer2_outputs(7099);
    outputs(7404) <= not(layer2_outputs(1256));
    outputs(7405) <= not((layer2_outputs(9256)) xor (layer2_outputs(7342)));
    outputs(7406) <= not(layer2_outputs(9822));
    outputs(7407) <= not((layer2_outputs(1030)) xor (layer2_outputs(10206)));
    outputs(7408) <= not((layer2_outputs(516)) or (layer2_outputs(2501)));
    outputs(7409) <= not((layer2_outputs(1293)) xor (layer2_outputs(9030)));
    outputs(7410) <= not(layer2_outputs(5903));
    outputs(7411) <= layer2_outputs(9215);
    outputs(7412) <= layer2_outputs(2216);
    outputs(7413) <= not((layer2_outputs(9913)) and (layer2_outputs(9652)));
    outputs(7414) <= (layer2_outputs(5782)) xor (layer2_outputs(6566));
    outputs(7415) <= not(layer2_outputs(9326));
    outputs(7416) <= not((layer2_outputs(7411)) or (layer2_outputs(3420)));
    outputs(7417) <= (layer2_outputs(415)) and not (layer2_outputs(6829));
    outputs(7418) <= not(layer2_outputs(3533));
    outputs(7419) <= (layer2_outputs(2586)) xor (layer2_outputs(4889));
    outputs(7420) <= layer2_outputs(9179);
    outputs(7421) <= not(layer2_outputs(8732));
    outputs(7422) <= layer2_outputs(2767);
    outputs(7423) <= not((layer2_outputs(8988)) xor (layer2_outputs(8134)));
    outputs(7424) <= (layer2_outputs(1949)) and (layer2_outputs(7885));
    outputs(7425) <= layer2_outputs(10038);
    outputs(7426) <= not(layer2_outputs(4990));
    outputs(7427) <= (layer2_outputs(6497)) and not (layer2_outputs(9707));
    outputs(7428) <= not((layer2_outputs(5695)) or (layer2_outputs(3475)));
    outputs(7429) <= not(layer2_outputs(1856));
    outputs(7430) <= (layer2_outputs(2540)) and not (layer2_outputs(2955));
    outputs(7431) <= layer2_outputs(2051);
    outputs(7432) <= not((layer2_outputs(3777)) xor (layer2_outputs(8406)));
    outputs(7433) <= (layer2_outputs(2814)) and (layer2_outputs(2971));
    outputs(7434) <= not((layer2_outputs(4137)) xor (layer2_outputs(1579)));
    outputs(7435) <= not(layer2_outputs(4820));
    outputs(7436) <= (layer2_outputs(4456)) xor (layer2_outputs(4781));
    outputs(7437) <= not(layer2_outputs(6786));
    outputs(7438) <= not((layer2_outputs(417)) xor (layer2_outputs(9407)));
    outputs(7439) <= not(layer2_outputs(1338));
    outputs(7440) <= not((layer2_outputs(9886)) xor (layer2_outputs(7400)));
    outputs(7441) <= (layer2_outputs(5808)) and not (layer2_outputs(435));
    outputs(7442) <= not((layer2_outputs(10217)) xor (layer2_outputs(9162)));
    outputs(7443) <= not(layer2_outputs(3238));
    outputs(7444) <= (layer2_outputs(2644)) xor (layer2_outputs(1272));
    outputs(7445) <= not((layer2_outputs(5131)) xor (layer2_outputs(8839)));
    outputs(7446) <= (layer2_outputs(9848)) and not (layer2_outputs(6321));
    outputs(7447) <= not(layer2_outputs(1220));
    outputs(7448) <= (layer2_outputs(8575)) xor (layer2_outputs(4995));
    outputs(7449) <= not((layer2_outputs(750)) xor (layer2_outputs(1345)));
    outputs(7450) <= (layer2_outputs(3470)) xor (layer2_outputs(7983));
    outputs(7451) <= (layer2_outputs(7705)) xor (layer2_outputs(7161));
    outputs(7452) <= not(layer2_outputs(3479));
    outputs(7453) <= layer2_outputs(5479);
    outputs(7454) <= layer2_outputs(3496);
    outputs(7455) <= layer2_outputs(5644);
    outputs(7456) <= (layer2_outputs(3373)) or (layer2_outputs(4336));
    outputs(7457) <= not((layer2_outputs(4436)) xor (layer2_outputs(3841)));
    outputs(7458) <= layer2_outputs(2268);
    outputs(7459) <= (layer2_outputs(9113)) and not (layer2_outputs(5460));
    outputs(7460) <= (layer2_outputs(9940)) and not (layer2_outputs(5705));
    outputs(7461) <= not((layer2_outputs(9539)) xor (layer2_outputs(5974)));
    outputs(7462) <= layer2_outputs(4022);
    outputs(7463) <= not((layer2_outputs(2185)) xor (layer2_outputs(261)));
    outputs(7464) <= not(layer2_outputs(3392));
    outputs(7465) <= layer2_outputs(10047);
    outputs(7466) <= (layer2_outputs(3536)) and (layer2_outputs(7020));
    outputs(7467) <= layer2_outputs(2172);
    outputs(7468) <= layer2_outputs(3698);
    outputs(7469) <= not(layer2_outputs(915));
    outputs(7470) <= not(layer2_outputs(5319));
    outputs(7471) <= layer2_outputs(2290);
    outputs(7472) <= not(layer2_outputs(4859));
    outputs(7473) <= not(layer2_outputs(3097));
    outputs(7474) <= not((layer2_outputs(5825)) xor (layer2_outputs(2242)));
    outputs(7475) <= layer2_outputs(3071);
    outputs(7476) <= not(layer2_outputs(2034));
    outputs(7477) <= not(layer2_outputs(10098)) or (layer2_outputs(2215));
    outputs(7478) <= not(layer2_outputs(8066));
    outputs(7479) <= (layer2_outputs(2216)) and (layer2_outputs(6269));
    outputs(7480) <= not(layer2_outputs(4133));
    outputs(7481) <= (layer2_outputs(10111)) and not (layer2_outputs(7565));
    outputs(7482) <= not((layer2_outputs(7275)) and (layer2_outputs(791)));
    outputs(7483) <= not(layer2_outputs(2813));
    outputs(7484) <= layer2_outputs(107);
    outputs(7485) <= not(layer2_outputs(269));
    outputs(7486) <= (layer2_outputs(8456)) and (layer2_outputs(2904));
    outputs(7487) <= layer2_outputs(9525);
    outputs(7488) <= (layer2_outputs(1298)) xor (layer2_outputs(408));
    outputs(7489) <= not((layer2_outputs(6741)) and (layer2_outputs(9301)));
    outputs(7490) <= not(layer2_outputs(7875));
    outputs(7491) <= layer2_outputs(1409);
    outputs(7492) <= (layer2_outputs(4250)) and not (layer2_outputs(6822));
    outputs(7493) <= layer2_outputs(10164);
    outputs(7494) <= not(layer2_outputs(8973));
    outputs(7495) <= not(layer2_outputs(7470)) or (layer2_outputs(129));
    outputs(7496) <= not((layer2_outputs(6030)) xor (layer2_outputs(3346)));
    outputs(7497) <= layer2_outputs(1051);
    outputs(7498) <= not(layer2_outputs(2054));
    outputs(7499) <= layer2_outputs(6570);
    outputs(7500) <= (layer2_outputs(4409)) xor (layer2_outputs(2467));
    outputs(7501) <= not(layer2_outputs(10120));
    outputs(7502) <= layer2_outputs(5430);
    outputs(7503) <= not((layer2_outputs(5162)) and (layer2_outputs(6145)));
    outputs(7504) <= not((layer2_outputs(9162)) or (layer2_outputs(7434)));
    outputs(7505) <= layer2_outputs(8375);
    outputs(7506) <= not(layer2_outputs(9337));
    outputs(7507) <= not((layer2_outputs(8568)) xor (layer2_outputs(9054)));
    outputs(7508) <= not((layer2_outputs(1112)) xor (layer2_outputs(7405)));
    outputs(7509) <= (layer2_outputs(7131)) and not (layer2_outputs(2009));
    outputs(7510) <= layer2_outputs(10127);
    outputs(7511) <= layer2_outputs(7374);
    outputs(7512) <= layer2_outputs(7728);
    outputs(7513) <= layer2_outputs(6578);
    outputs(7514) <= not((layer2_outputs(1947)) or (layer2_outputs(2968)));
    outputs(7515) <= not(layer2_outputs(1672));
    outputs(7516) <= not(layer2_outputs(8105));
    outputs(7517) <= layer2_outputs(7454);
    outputs(7518) <= not(layer2_outputs(3614));
    outputs(7519) <= not((layer2_outputs(1860)) xor (layer2_outputs(5553)));
    outputs(7520) <= layer2_outputs(7250);
    outputs(7521) <= not(layer2_outputs(6235));
    outputs(7522) <= layer2_outputs(9703);
    outputs(7523) <= (layer2_outputs(6737)) and not (layer2_outputs(1510));
    outputs(7524) <= not(layer2_outputs(5104));
    outputs(7525) <= (layer2_outputs(2953)) xor (layer2_outputs(1996));
    outputs(7526) <= (layer2_outputs(21)) xor (layer2_outputs(7449));
    outputs(7527) <= layer2_outputs(5832);
    outputs(7528) <= (layer2_outputs(271)) or (layer2_outputs(2560));
    outputs(7529) <= not(layer2_outputs(206));
    outputs(7530) <= not(layer2_outputs(5360));
    outputs(7531) <= not((layer2_outputs(3275)) xor (layer2_outputs(8865)));
    outputs(7532) <= not(layer2_outputs(7706));
    outputs(7533) <= (layer2_outputs(3068)) or (layer2_outputs(3252));
    outputs(7534) <= (layer2_outputs(9700)) and not (layer2_outputs(9642));
    outputs(7535) <= not(layer2_outputs(644));
    outputs(7536) <= layer2_outputs(9340);
    outputs(7537) <= (layer2_outputs(5585)) and not (layer2_outputs(9078));
    outputs(7538) <= not((layer2_outputs(7131)) xor (layer2_outputs(5446)));
    outputs(7539) <= (layer2_outputs(5249)) and not (layer2_outputs(9654));
    outputs(7540) <= (layer2_outputs(4148)) and not (layer2_outputs(3895));
    outputs(7541) <= not(layer2_outputs(156));
    outputs(7542) <= (layer2_outputs(8899)) and (layer2_outputs(9149));
    outputs(7543) <= not(layer2_outputs(5362));
    outputs(7544) <= not(layer2_outputs(1403));
    outputs(7545) <= layer2_outputs(6116);
    outputs(7546) <= not(layer2_outputs(1153));
    outputs(7547) <= layer2_outputs(820);
    outputs(7548) <= (layer2_outputs(368)) xor (layer2_outputs(493));
    outputs(7549) <= layer2_outputs(5038);
    outputs(7550) <= not((layer2_outputs(5864)) xor (layer2_outputs(829)));
    outputs(7551) <= not(layer2_outputs(7975));
    outputs(7552) <= (layer2_outputs(9238)) and not (layer2_outputs(10218));
    outputs(7553) <= (layer2_outputs(397)) and not (layer2_outputs(1021));
    outputs(7554) <= not(layer2_outputs(5790));
    outputs(7555) <= not(layer2_outputs(1554));
    outputs(7556) <= not(layer2_outputs(6584));
    outputs(7557) <= layer2_outputs(7704);
    outputs(7558) <= (layer2_outputs(8295)) and (layer2_outputs(5684));
    outputs(7559) <= (layer2_outputs(3919)) xor (layer2_outputs(1147));
    outputs(7560) <= not(layer2_outputs(2038)) or (layer2_outputs(1218));
    outputs(7561) <= (layer2_outputs(8937)) xor (layer2_outputs(3503));
    outputs(7562) <= not(layer2_outputs(602));
    outputs(7563) <= layer2_outputs(2183);
    outputs(7564) <= layer2_outputs(7843);
    outputs(7565) <= (layer2_outputs(1017)) xor (layer2_outputs(8870));
    outputs(7566) <= not((layer2_outputs(9900)) xor (layer2_outputs(477)));
    outputs(7567) <= layer2_outputs(5758);
    outputs(7568) <= layer2_outputs(1158);
    outputs(7569) <= not(layer2_outputs(9982));
    outputs(7570) <= not(layer2_outputs(1306)) or (layer2_outputs(5972));
    outputs(7571) <= not((layer2_outputs(9373)) or (layer2_outputs(5741)));
    outputs(7572) <= (layer2_outputs(7022)) and (layer2_outputs(2423));
    outputs(7573) <= not((layer2_outputs(918)) xor (layer2_outputs(356)));
    outputs(7574) <= not(layer2_outputs(4878));
    outputs(7575) <= (layer2_outputs(6590)) xor (layer2_outputs(495));
    outputs(7576) <= (layer2_outputs(9362)) and not (layer2_outputs(9043));
    outputs(7577) <= layer2_outputs(6299);
    outputs(7578) <= layer2_outputs(221);
    outputs(7579) <= not((layer2_outputs(466)) xor (layer2_outputs(8300)));
    outputs(7580) <= (layer2_outputs(9624)) xor (layer2_outputs(3808));
    outputs(7581) <= not((layer2_outputs(8594)) xor (layer2_outputs(9816)));
    outputs(7582) <= layer2_outputs(1714);
    outputs(7583) <= layer2_outputs(9055);
    outputs(7584) <= layer2_outputs(8171);
    outputs(7585) <= (layer2_outputs(1212)) xor (layer2_outputs(2288));
    outputs(7586) <= (layer2_outputs(7643)) and not (layer2_outputs(9672));
    outputs(7587) <= (layer2_outputs(2983)) and not (layer2_outputs(6495));
    outputs(7588) <= layer2_outputs(1127);
    outputs(7589) <= layer2_outputs(10147);
    outputs(7590) <= (layer2_outputs(3801)) and not (layer2_outputs(9889));
    outputs(7591) <= layer2_outputs(274);
    outputs(7592) <= not((layer2_outputs(10130)) or (layer2_outputs(5027)));
    outputs(7593) <= not(layer2_outputs(8939));
    outputs(7594) <= layer2_outputs(2819);
    outputs(7595) <= not((layer2_outputs(7002)) xor (layer2_outputs(2219)));
    outputs(7596) <= not(layer2_outputs(8651));
    outputs(7597) <= not(layer2_outputs(5411));
    outputs(7598) <= layer2_outputs(6753);
    outputs(7599) <= layer2_outputs(747);
    outputs(7600) <= layer2_outputs(1966);
    outputs(7601) <= not(layer2_outputs(10104)) or (layer2_outputs(526));
    outputs(7602) <= layer2_outputs(2706);
    outputs(7603) <= not(layer2_outputs(5762));
    outputs(7604) <= layer2_outputs(2214);
    outputs(7605) <= layer2_outputs(3490);
    outputs(7606) <= layer2_outputs(9848);
    outputs(7607) <= not(layer2_outputs(1987));
    outputs(7608) <= not((layer2_outputs(6411)) or (layer2_outputs(6626)));
    outputs(7609) <= not(layer2_outputs(4086));
    outputs(7610) <= layer2_outputs(502);
    outputs(7611) <= not((layer2_outputs(8080)) xor (layer2_outputs(1382)));
    outputs(7612) <= layer2_outputs(9320);
    outputs(7613) <= not(layer2_outputs(6035));
    outputs(7614) <= (layer2_outputs(4884)) and not (layer2_outputs(10018));
    outputs(7615) <= (layer2_outputs(4288)) or (layer2_outputs(5893));
    outputs(7616) <= not((layer2_outputs(5492)) xor (layer2_outputs(6134)));
    outputs(7617) <= not(layer2_outputs(1761));
    outputs(7618) <= not((layer2_outputs(2906)) xor (layer2_outputs(8495)));
    outputs(7619) <= layer2_outputs(5712);
    outputs(7620) <= layer2_outputs(1089);
    outputs(7621) <= (layer2_outputs(9214)) and (layer2_outputs(2090));
    outputs(7622) <= (layer2_outputs(8242)) xor (layer2_outputs(2985));
    outputs(7623) <= not((layer2_outputs(9654)) xor (layer2_outputs(7913)));
    outputs(7624) <= layer2_outputs(9827);
    outputs(7625) <= layer2_outputs(4186);
    outputs(7626) <= not(layer2_outputs(6860));
    outputs(7627) <= layer2_outputs(3343);
    outputs(7628) <= (layer2_outputs(9414)) and not (layer2_outputs(7279));
    outputs(7629) <= not(layer2_outputs(3972));
    outputs(7630) <= layer2_outputs(9842);
    outputs(7631) <= (layer2_outputs(7238)) xor (layer2_outputs(1267));
    outputs(7632) <= not(layer2_outputs(5641));
    outputs(7633) <= not((layer2_outputs(7293)) xor (layer2_outputs(1956)));
    outputs(7634) <= not((layer2_outputs(5870)) xor (layer2_outputs(7897)));
    outputs(7635) <= (layer2_outputs(9400)) and not (layer2_outputs(10002));
    outputs(7636) <= not(layer2_outputs(3126));
    outputs(7637) <= not(layer2_outputs(4719));
    outputs(7638) <= not(layer2_outputs(8884));
    outputs(7639) <= (layer2_outputs(1606)) and (layer2_outputs(7590));
    outputs(7640) <= layer2_outputs(6443);
    outputs(7641) <= not(layer2_outputs(5679));
    outputs(7642) <= layer2_outputs(4632);
    outputs(7643) <= not(layer2_outputs(355));
    outputs(7644) <= layer2_outputs(9422);
    outputs(7645) <= layer2_outputs(7796);
    outputs(7646) <= layer2_outputs(873);
    outputs(7647) <= not((layer2_outputs(2972)) or (layer2_outputs(5120)));
    outputs(7648) <= not(layer2_outputs(1804));
    outputs(7649) <= layer2_outputs(2059);
    outputs(7650) <= not(layer2_outputs(3584)) or (layer2_outputs(5485));
    outputs(7651) <= (layer2_outputs(7164)) and not (layer2_outputs(10052));
    outputs(7652) <= layer2_outputs(5769);
    outputs(7653) <= layer2_outputs(4994);
    outputs(7654) <= (layer2_outputs(8064)) and (layer2_outputs(3112));
    outputs(7655) <= not(layer2_outputs(1251));
    outputs(7656) <= not((layer2_outputs(704)) or (layer2_outputs(9191)));
    outputs(7657) <= (layer2_outputs(4967)) and not (layer2_outputs(4246));
    outputs(7658) <= layer2_outputs(2673);
    outputs(7659) <= (layer2_outputs(8955)) xor (layer2_outputs(1543));
    outputs(7660) <= not(layer2_outputs(1811));
    outputs(7661) <= layer2_outputs(3562);
    outputs(7662) <= not(layer2_outputs(3905));
    outputs(7663) <= layer2_outputs(9045);
    outputs(7664) <= (layer2_outputs(4023)) and not (layer2_outputs(2526));
    outputs(7665) <= layer2_outputs(7325);
    outputs(7666) <= not(layer2_outputs(3685));
    outputs(7667) <= not(layer2_outputs(6879));
    outputs(7668) <= (layer2_outputs(485)) or (layer2_outputs(8411));
    outputs(7669) <= not(layer2_outputs(1008));
    outputs(7670) <= not(layer2_outputs(8964));
    outputs(7671) <= not(layer2_outputs(10060));
    outputs(7672) <= layer2_outputs(7330);
    outputs(7673) <= not(layer2_outputs(9303));
    outputs(7674) <= (layer2_outputs(9995)) xor (layer2_outputs(909));
    outputs(7675) <= not(layer2_outputs(5504));
    outputs(7676) <= layer2_outputs(9418);
    outputs(7677) <= not(layer2_outputs(3255));
    outputs(7678) <= layer2_outputs(742);
    outputs(7679) <= (layer2_outputs(475)) and not (layer2_outputs(4711));
    outputs(7680) <= not(layer2_outputs(2669));
    outputs(7681) <= not(layer2_outputs(1320));
    outputs(7682) <= (layer2_outputs(8126)) xor (layer2_outputs(7929));
    outputs(7683) <= (layer2_outputs(10037)) and not (layer2_outputs(7203));
    outputs(7684) <= not(layer2_outputs(3100)) or (layer2_outputs(1666));
    outputs(7685) <= not(layer2_outputs(6700));
    outputs(7686) <= (layer2_outputs(8329)) and not (layer2_outputs(833));
    outputs(7687) <= not((layer2_outputs(1798)) xor (layer2_outputs(2021)));
    outputs(7688) <= layer2_outputs(9006);
    outputs(7689) <= not((layer2_outputs(2077)) xor (layer2_outputs(2501)));
    outputs(7690) <= (layer2_outputs(1021)) xor (layer2_outputs(948));
    outputs(7691) <= layer2_outputs(9657);
    outputs(7692) <= layer2_outputs(7795);
    outputs(7693) <= not(layer2_outputs(7710));
    outputs(7694) <= not(layer2_outputs(4584));
    outputs(7695) <= (layer2_outputs(3477)) and not (layer2_outputs(427));
    outputs(7696) <= layer2_outputs(2361);
    outputs(7697) <= not((layer2_outputs(4599)) xor (layer2_outputs(216)));
    outputs(7698) <= (layer2_outputs(7891)) xor (layer2_outputs(1877));
    outputs(7699) <= layer2_outputs(9926);
    outputs(7700) <= layer2_outputs(6890);
    outputs(7701) <= not(layer2_outputs(1333));
    outputs(7702) <= not(layer2_outputs(4360));
    outputs(7703) <= not((layer2_outputs(7727)) xor (layer2_outputs(1788)));
    outputs(7704) <= layer2_outputs(6753);
    outputs(7705) <= (layer2_outputs(5857)) and not (layer2_outputs(839));
    outputs(7706) <= not(layer2_outputs(504));
    outputs(7707) <= layer2_outputs(3753);
    outputs(7708) <= not(layer2_outputs(9599));
    outputs(7709) <= not((layer2_outputs(8689)) xor (layer2_outputs(2221)));
    outputs(7710) <= not((layer2_outputs(7735)) xor (layer2_outputs(7816)));
    outputs(7711) <= (layer2_outputs(2866)) xor (layer2_outputs(2660));
    outputs(7712) <= layer2_outputs(6176);
    outputs(7713) <= layer2_outputs(4618);
    outputs(7714) <= not((layer2_outputs(1810)) xor (layer2_outputs(8971)));
    outputs(7715) <= (layer2_outputs(9341)) and not (layer2_outputs(7560));
    outputs(7716) <= layer2_outputs(4389);
    outputs(7717) <= (layer2_outputs(5117)) and (layer2_outputs(8366));
    outputs(7718) <= layer2_outputs(8159);
    outputs(7719) <= layer2_outputs(10147);
    outputs(7720) <= not(layer2_outputs(2528));
    outputs(7721) <= not((layer2_outputs(6697)) xor (layer2_outputs(6190)));
    outputs(7722) <= (layer2_outputs(2870)) and not (layer2_outputs(4774));
    outputs(7723) <= layer2_outputs(1069);
    outputs(7724) <= layer2_outputs(6304);
    outputs(7725) <= not((layer2_outputs(1601)) xor (layer2_outputs(1100)));
    outputs(7726) <= not(layer2_outputs(7051));
    outputs(7727) <= not(layer2_outputs(5362));
    outputs(7728) <= layer2_outputs(9028);
    outputs(7729) <= not(layer2_outputs(2548));
    outputs(7730) <= (layer2_outputs(4537)) and not (layer2_outputs(2149));
    outputs(7731) <= not(layer2_outputs(6799)) or (layer2_outputs(3425));
    outputs(7732) <= not(layer2_outputs(5982));
    outputs(7733) <= not((layer2_outputs(7355)) xor (layer2_outputs(1067)));
    outputs(7734) <= not((layer2_outputs(6075)) xor (layer2_outputs(5095)));
    outputs(7735) <= layer2_outputs(4883);
    outputs(7736) <= layer2_outputs(3873);
    outputs(7737) <= (layer2_outputs(3689)) and not (layer2_outputs(1336));
    outputs(7738) <= layer2_outputs(4199);
    outputs(7739) <= not(layer2_outputs(7481));
    outputs(7740) <= (layer2_outputs(7080)) xor (layer2_outputs(7466));
    outputs(7741) <= (layer2_outputs(2805)) and not (layer2_outputs(7223));
    outputs(7742) <= layer2_outputs(3035);
    outputs(7743) <= not((layer2_outputs(2723)) xor (layer2_outputs(5136)));
    outputs(7744) <= layer2_outputs(5832);
    outputs(7745) <= layer2_outputs(7099);
    outputs(7746) <= layer2_outputs(8557);
    outputs(7747) <= layer2_outputs(2774);
    outputs(7748) <= not((layer2_outputs(2394)) xor (layer2_outputs(6915)));
    outputs(7749) <= not((layer2_outputs(8857)) xor (layer2_outputs(6492)));
    outputs(7750) <= (layer2_outputs(3167)) and not (layer2_outputs(3475));
    outputs(7751) <= (layer2_outputs(6125)) or (layer2_outputs(160));
    outputs(7752) <= not(layer2_outputs(933));
    outputs(7753) <= not(layer2_outputs(1716));
    outputs(7754) <= (layer2_outputs(7778)) and not (layer2_outputs(7237));
    outputs(7755) <= not((layer2_outputs(1335)) xor (layer2_outputs(259)));
    outputs(7756) <= not(layer2_outputs(7634));
    outputs(7757) <= (layer2_outputs(9064)) xor (layer2_outputs(3546));
    outputs(7758) <= (layer2_outputs(5465)) and not (layer2_outputs(6786));
    outputs(7759) <= (layer2_outputs(8015)) and not (layer2_outputs(9457));
    outputs(7760) <= not(layer2_outputs(3951));
    outputs(7761) <= not(layer2_outputs(4433));
    outputs(7762) <= not((layer2_outputs(2452)) xor (layer2_outputs(9077)));
    outputs(7763) <= layer2_outputs(4280);
    outputs(7764) <= layer2_outputs(4447);
    outputs(7765) <= not((layer2_outputs(1580)) or (layer2_outputs(1002)));
    outputs(7766) <= not(layer2_outputs(3837));
    outputs(7767) <= not((layer2_outputs(3293)) xor (layer2_outputs(4585)));
    outputs(7768) <= layer2_outputs(499);
    outputs(7769) <= not(layer2_outputs(6267));
    outputs(7770) <= not(layer2_outputs(8590));
    outputs(7771) <= not(layer2_outputs(3063));
    outputs(7772) <= layer2_outputs(6338);
    outputs(7773) <= layer2_outputs(468);
    outputs(7774) <= layer2_outputs(5807);
    outputs(7775) <= (layer2_outputs(10162)) and not (layer2_outputs(3652));
    outputs(7776) <= layer2_outputs(7912);
    outputs(7777) <= layer2_outputs(276);
    outputs(7778) <= (layer2_outputs(6136)) and not (layer2_outputs(5250));
    outputs(7779) <= (layer2_outputs(7186)) xor (layer2_outputs(5780));
    outputs(7780) <= layer2_outputs(7030);
    outputs(7781) <= not((layer2_outputs(3483)) xor (layer2_outputs(2086)));
    outputs(7782) <= (layer2_outputs(1083)) and not (layer2_outputs(696));
    outputs(7783) <= (layer2_outputs(9846)) xor (layer2_outputs(5715));
    outputs(7784) <= not(layer2_outputs(4820));
    outputs(7785) <= (layer2_outputs(5609)) xor (layer2_outputs(10163));
    outputs(7786) <= layer2_outputs(1959);
    outputs(7787) <= not(layer2_outputs(94));
    outputs(7788) <= not(layer2_outputs(8719));
    outputs(7789) <= (layer2_outputs(5289)) xor (layer2_outputs(6599));
    outputs(7790) <= (layer2_outputs(7501)) xor (layer2_outputs(1797));
    outputs(7791) <= not((layer2_outputs(3132)) or (layer2_outputs(1602)));
    outputs(7792) <= layer2_outputs(9602);
    outputs(7793) <= not(layer2_outputs(9825));
    outputs(7794) <= (layer2_outputs(4363)) xor (layer2_outputs(7270));
    outputs(7795) <= not(layer2_outputs(4160));
    outputs(7796) <= not((layer2_outputs(331)) and (layer2_outputs(4370)));
    outputs(7797) <= layer2_outputs(2050);
    outputs(7798) <= not(layer2_outputs(8030));
    outputs(7799) <= layer2_outputs(8407);
    outputs(7800) <= not(layer2_outputs(9872));
    outputs(7801) <= not(layer2_outputs(7256));
    outputs(7802) <= (layer2_outputs(7925)) xor (layer2_outputs(1057));
    outputs(7803) <= layer2_outputs(4116);
    outputs(7804) <= (layer2_outputs(8151)) and not (layer2_outputs(2016));
    outputs(7805) <= not((layer2_outputs(8784)) or (layer2_outputs(5996)));
    outputs(7806) <= layer2_outputs(3001);
    outputs(7807) <= (layer2_outputs(8367)) and not (layer2_outputs(5358));
    outputs(7808) <= layer2_outputs(1574);
    outputs(7809) <= (layer2_outputs(474)) and (layer2_outputs(3859));
    outputs(7810) <= (layer2_outputs(966)) and not (layer2_outputs(5183));
    outputs(7811) <= not((layer2_outputs(279)) or (layer2_outputs(7601)));
    outputs(7812) <= layer2_outputs(8511);
    outputs(7813) <= not(layer2_outputs(4603));
    outputs(7814) <= not(layer2_outputs(7051));
    outputs(7815) <= layer2_outputs(539);
    outputs(7816) <= layer2_outputs(10069);
    outputs(7817) <= layer2_outputs(7192);
    outputs(7818) <= layer2_outputs(6496);
    outputs(7819) <= not(layer2_outputs(9804));
    outputs(7820) <= not(layer2_outputs(3135));
    outputs(7821) <= not(layer2_outputs(4996));
    outputs(7822) <= layer2_outputs(201);
    outputs(7823) <= not(layer2_outputs(6383));
    outputs(7824) <= (layer2_outputs(1422)) and (layer2_outputs(5484));
    outputs(7825) <= not(layer2_outputs(8828));
    outputs(7826) <= not(layer2_outputs(222)) or (layer2_outputs(3300));
    outputs(7827) <= layer2_outputs(5024);
    outputs(7828) <= layer2_outputs(4321);
    outputs(7829) <= not(layer2_outputs(9402));
    outputs(7830) <= layer2_outputs(9283);
    outputs(7831) <= not(layer2_outputs(2973));
    outputs(7832) <= layer2_outputs(2339);
    outputs(7833) <= not(layer2_outputs(9268));
    outputs(7834) <= not((layer2_outputs(4579)) xor (layer2_outputs(1962)));
    outputs(7835) <= (layer2_outputs(5751)) xor (layer2_outputs(6506));
    outputs(7836) <= not((layer2_outputs(4597)) xor (layer2_outputs(2367)));
    outputs(7837) <= not(layer2_outputs(6986));
    outputs(7838) <= layer2_outputs(1148);
    outputs(7839) <= layer2_outputs(7555);
    outputs(7840) <= not(layer2_outputs(69));
    outputs(7841) <= layer2_outputs(3726);
    outputs(7842) <= layer2_outputs(7477);
    outputs(7843) <= layer2_outputs(9126);
    outputs(7844) <= not(layer2_outputs(6874));
    outputs(7845) <= not((layer2_outputs(9919)) xor (layer2_outputs(1152)));
    outputs(7846) <= not(layer2_outputs(9356)) or (layer2_outputs(4849));
    outputs(7847) <= not(layer2_outputs(3837));
    outputs(7848) <= (layer2_outputs(1525)) xor (layer2_outputs(6969));
    outputs(7849) <= layer2_outputs(3645);
    outputs(7850) <= layer2_outputs(8010);
    outputs(7851) <= layer2_outputs(1093);
    outputs(7852) <= (layer2_outputs(3524)) or (layer2_outputs(1201));
    outputs(7853) <= (layer2_outputs(1539)) xor (layer2_outputs(2411));
    outputs(7854) <= layer2_outputs(4897);
    outputs(7855) <= not((layer2_outputs(7048)) xor (layer2_outputs(6596)));
    outputs(7856) <= not((layer2_outputs(6503)) or (layer2_outputs(3123)));
    outputs(7857) <= layer2_outputs(3515);
    outputs(7858) <= layer2_outputs(8257);
    outputs(7859) <= (layer2_outputs(7266)) xor (layer2_outputs(6959));
    outputs(7860) <= not((layer2_outputs(5349)) xor (layer2_outputs(5283)));
    outputs(7861) <= not(layer2_outputs(1250));
    outputs(7862) <= (layer2_outputs(7417)) and not (layer2_outputs(6842));
    outputs(7863) <= (layer2_outputs(3066)) and not (layer2_outputs(6221));
    outputs(7864) <= not(layer2_outputs(8945));
    outputs(7865) <= layer2_outputs(8835);
    outputs(7866) <= not(layer2_outputs(7111));
    outputs(7867) <= not(layer2_outputs(8589));
    outputs(7868) <= not(layer2_outputs(5838));
    outputs(7869) <= (layer2_outputs(9699)) and not (layer2_outputs(1579));
    outputs(7870) <= layer2_outputs(5582);
    outputs(7871) <= not((layer2_outputs(3357)) xor (layer2_outputs(2328)));
    outputs(7872) <= not(layer2_outputs(9959));
    outputs(7873) <= layer2_outputs(629);
    outputs(7874) <= (layer2_outputs(117)) xor (layer2_outputs(5969));
    outputs(7875) <= not((layer2_outputs(9577)) or (layer2_outputs(4842)));
    outputs(7876) <= layer2_outputs(4249);
    outputs(7877) <= layer2_outputs(1587);
    outputs(7878) <= layer2_outputs(2378);
    outputs(7879) <= not(layer2_outputs(258));
    outputs(7880) <= layer2_outputs(8181);
    outputs(7881) <= (layer2_outputs(8477)) xor (layer2_outputs(830));
    outputs(7882) <= (layer2_outputs(7074)) xor (layer2_outputs(3079));
    outputs(7883) <= layer2_outputs(8605);
    outputs(7884) <= (layer2_outputs(8091)) and (layer2_outputs(9678));
    outputs(7885) <= not(layer2_outputs(6553));
    outputs(7886) <= not(layer2_outputs(1284));
    outputs(7887) <= (layer2_outputs(4740)) and not (layer2_outputs(2156));
    outputs(7888) <= layer2_outputs(2814);
    outputs(7889) <= not(layer2_outputs(3601));
    outputs(7890) <= layer2_outputs(4986);
    outputs(7891) <= not(layer2_outputs(6899));
    outputs(7892) <= layer2_outputs(5102);
    outputs(7893) <= layer2_outputs(3593);
    outputs(7894) <= not(layer2_outputs(4211));
    outputs(7895) <= not(layer2_outputs(3738));
    outputs(7896) <= layer2_outputs(3554);
    outputs(7897) <= not(layer2_outputs(1898));
    outputs(7898) <= not(layer2_outputs(5457));
    outputs(7899) <= (layer2_outputs(10131)) xor (layer2_outputs(3016));
    outputs(7900) <= (layer2_outputs(7566)) and (layer2_outputs(4906));
    outputs(7901) <= (layer2_outputs(8528)) and (layer2_outputs(3124));
    outputs(7902) <= not(layer2_outputs(8928));
    outputs(7903) <= (layer2_outputs(1217)) and not (layer2_outputs(3415));
    outputs(7904) <= layer2_outputs(4525);
    outputs(7905) <= not((layer2_outputs(1144)) and (layer2_outputs(6597)));
    outputs(7906) <= layer2_outputs(8888);
    outputs(7907) <= not(layer2_outputs(6894));
    outputs(7908) <= layer2_outputs(2260);
    outputs(7909) <= layer2_outputs(2954);
    outputs(7910) <= (layer2_outputs(3933)) xor (layer2_outputs(7856));
    outputs(7911) <= not(layer2_outputs(4812)) or (layer2_outputs(1329));
    outputs(7912) <= layer2_outputs(2430);
    outputs(7913) <= not(layer2_outputs(264)) or (layer2_outputs(8624));
    outputs(7914) <= not((layer2_outputs(3354)) xor (layer2_outputs(4898)));
    outputs(7915) <= (layer2_outputs(7519)) and not (layer2_outputs(8637));
    outputs(7916) <= (layer2_outputs(3021)) and (layer2_outputs(9246));
    outputs(7917) <= not(layer2_outputs(959));
    outputs(7918) <= layer2_outputs(5781);
    outputs(7919) <= (layer2_outputs(2314)) xor (layer2_outputs(12));
    outputs(7920) <= layer2_outputs(3281);
    outputs(7921) <= not(layer2_outputs(4134));
    outputs(7922) <= not(layer2_outputs(5551)) or (layer2_outputs(655));
    outputs(7923) <= layer2_outputs(6771);
    outputs(7924) <= layer2_outputs(8980);
    outputs(7925) <= not(layer2_outputs(4859));
    outputs(7926) <= not(layer2_outputs(4530));
    outputs(7927) <= not(layer2_outputs(5355));
    outputs(7928) <= (layer2_outputs(2034)) xor (layer2_outputs(7400));
    outputs(7929) <= (layer2_outputs(7393)) and (layer2_outputs(4272));
    outputs(7930) <= (layer2_outputs(3090)) and not (layer2_outputs(1598));
    outputs(7931) <= (layer2_outputs(4300)) and not (layer2_outputs(7106));
    outputs(7932) <= not((layer2_outputs(3062)) xor (layer2_outputs(797)));
    outputs(7933) <= (layer2_outputs(3389)) xor (layer2_outputs(5151));
    outputs(7934) <= (layer2_outputs(2753)) and not (layer2_outputs(9616));
    outputs(7935) <= (layer2_outputs(4616)) xor (layer2_outputs(7971));
    outputs(7936) <= (layer2_outputs(177)) and not (layer2_outputs(1604));
    outputs(7937) <= (layer2_outputs(5276)) xor (layer2_outputs(6421));
    outputs(7938) <= not(layer2_outputs(4710));
    outputs(7939) <= (layer2_outputs(8298)) and (layer2_outputs(6366));
    outputs(7940) <= not((layer2_outputs(1642)) or (layer2_outputs(8452)));
    outputs(7941) <= layer2_outputs(5542);
    outputs(7942) <= layer2_outputs(2210);
    outputs(7943) <= not(layer2_outputs(7004));
    outputs(7944) <= not(layer2_outputs(2177));
    outputs(7945) <= not(layer2_outputs(6969));
    outputs(7946) <= (layer2_outputs(7611)) xor (layer2_outputs(1866));
    outputs(7947) <= not(layer2_outputs(5070));
    outputs(7948) <= not((layer2_outputs(4452)) xor (layer2_outputs(7075)));
    outputs(7949) <= layer2_outputs(8381);
    outputs(7950) <= not(layer2_outputs(6380));
    outputs(7951) <= not(layer2_outputs(2264));
    outputs(7952) <= not((layer2_outputs(6433)) xor (layer2_outputs(2212)));
    outputs(7953) <= not(layer2_outputs(8945));
    outputs(7954) <= not(layer2_outputs(1517));
    outputs(7955) <= layer2_outputs(5773);
    outputs(7956) <= (layer2_outputs(3990)) and not (layer2_outputs(7823));
    outputs(7957) <= layer2_outputs(8614);
    outputs(7958) <= not((layer2_outputs(4893)) xor (layer2_outputs(9819)));
    outputs(7959) <= (layer2_outputs(324)) or (layer2_outputs(3308));
    outputs(7960) <= (layer2_outputs(6513)) and not (layer2_outputs(5777));
    outputs(7961) <= layer2_outputs(4808);
    outputs(7962) <= not(layer2_outputs(9696));
    outputs(7963) <= not(layer2_outputs(2289));
    outputs(7964) <= layer2_outputs(8987);
    outputs(7965) <= not(layer2_outputs(3291));
    outputs(7966) <= not((layer2_outputs(3298)) xor (layer2_outputs(2641)));
    outputs(7967) <= layer2_outputs(5028);
    outputs(7968) <= layer2_outputs(4188);
    outputs(7969) <= layer2_outputs(5113);
    outputs(7970) <= not((layer2_outputs(4550)) xor (layer2_outputs(6213)));
    outputs(7971) <= layer2_outputs(2799);
    outputs(7972) <= not(layer2_outputs(8110));
    outputs(7973) <= not((layer2_outputs(3813)) xor (layer2_outputs(6307)));
    outputs(7974) <= not(layer2_outputs(1398));
    outputs(7975) <= (layer2_outputs(709)) and not (layer2_outputs(665));
    outputs(7976) <= not((layer2_outputs(3081)) or (layer2_outputs(5468)));
    outputs(7977) <= not(layer2_outputs(1907));
    outputs(7978) <= layer2_outputs(4412);
    outputs(7979) <= (layer2_outputs(2136)) xor (layer2_outputs(9300));
    outputs(7980) <= layer2_outputs(6688);
    outputs(7981) <= not(layer2_outputs(3664));
    outputs(7982) <= not(layer2_outputs(2652));
    outputs(7983) <= layer2_outputs(4790);
    outputs(7984) <= not((layer2_outputs(4298)) and (layer2_outputs(7542)));
    outputs(7985) <= layer2_outputs(3040);
    outputs(7986) <= layer2_outputs(7293);
    outputs(7987) <= (layer2_outputs(8011)) and (layer2_outputs(7215));
    outputs(7988) <= (layer2_outputs(6127)) and not (layer2_outputs(9610));
    outputs(7989) <= not(layer2_outputs(615));
    outputs(7990) <= (layer2_outputs(9577)) xor (layer2_outputs(1317));
    outputs(7991) <= (layer2_outputs(6660)) and not (layer2_outputs(6000));
    outputs(7992) <= not((layer2_outputs(6917)) xor (layer2_outputs(9066)));
    outputs(7993) <= layer2_outputs(3322);
    outputs(7994) <= layer2_outputs(6932);
    outputs(7995) <= not((layer2_outputs(2951)) and (layer2_outputs(6149)));
    outputs(7996) <= not(layer2_outputs(472));
    outputs(7997) <= not((layer2_outputs(5944)) or (layer2_outputs(10224)));
    outputs(7998) <= not((layer2_outputs(9074)) xor (layer2_outputs(2434)));
    outputs(7999) <= layer2_outputs(8763);
    outputs(8000) <= not(layer2_outputs(8917));
    outputs(8001) <= layer2_outputs(9656);
    outputs(8002) <= not(layer2_outputs(8537));
    outputs(8003) <= (layer2_outputs(8152)) xor (layer2_outputs(1477));
    outputs(8004) <= layer2_outputs(4330);
    outputs(8005) <= not((layer2_outputs(4313)) or (layer2_outputs(8878)));
    outputs(8006) <= layer2_outputs(1344);
    outputs(8007) <= not(layer2_outputs(4067));
    outputs(8008) <= not(layer2_outputs(6781));
    outputs(8009) <= (layer2_outputs(6928)) and not (layer2_outputs(3173));
    outputs(8010) <= layer2_outputs(5884);
    outputs(8011) <= (layer2_outputs(7957)) xor (layer2_outputs(4900));
    outputs(8012) <= not((layer2_outputs(6752)) xor (layer2_outputs(6731)));
    outputs(8013) <= layer2_outputs(7888);
    outputs(8014) <= not(layer2_outputs(6437));
    outputs(8015) <= not(layer2_outputs(6178)) or (layer2_outputs(9095));
    outputs(8016) <= layer2_outputs(2015);
    outputs(8017) <= (layer2_outputs(182)) xor (layer2_outputs(8300));
    outputs(8018) <= layer2_outputs(6693);
    outputs(8019) <= not(layer2_outputs(455));
    outputs(8020) <= not(layer2_outputs(3355));
    outputs(8021) <= layer2_outputs(8851);
    outputs(8022) <= not(layer2_outputs(8658));
    outputs(8023) <= not(layer2_outputs(9339));
    outputs(8024) <= not(layer2_outputs(9606));
    outputs(8025) <= (layer2_outputs(2563)) or (layer2_outputs(9417));
    outputs(8026) <= layer2_outputs(8309);
    outputs(8027) <= not(layer2_outputs(2464));
    outputs(8028) <= not(layer2_outputs(2634));
    outputs(8029) <= layer2_outputs(2183);
    outputs(8030) <= (layer2_outputs(8347)) and (layer2_outputs(7642));
    outputs(8031) <= not((layer2_outputs(3761)) xor (layer2_outputs(6805)));
    outputs(8032) <= layer2_outputs(5907);
    outputs(8033) <= layer2_outputs(4973);
    outputs(8034) <= not((layer2_outputs(2745)) xor (layer2_outputs(856)));
    outputs(8035) <= layer2_outputs(1358);
    outputs(8036) <= layer2_outputs(6843);
    outputs(8037) <= layer2_outputs(9954);
    outputs(8038) <= (layer2_outputs(3712)) and not (layer2_outputs(6235));
    outputs(8039) <= (layer2_outputs(4390)) and (layer2_outputs(810));
    outputs(8040) <= layer2_outputs(4492);
    outputs(8041) <= layer2_outputs(3794);
    outputs(8042) <= not(layer2_outputs(6474));
    outputs(8043) <= not(layer2_outputs(1679));
    outputs(8044) <= (layer2_outputs(5501)) xor (layer2_outputs(6402));
    outputs(8045) <= layer2_outputs(7152);
    outputs(8046) <= layer2_outputs(7790);
    outputs(8047) <= layer2_outputs(9507);
    outputs(8048) <= not(layer2_outputs(8930));
    outputs(8049) <= layer2_outputs(3423);
    outputs(8050) <= (layer2_outputs(6639)) xor (layer2_outputs(7221));
    outputs(8051) <= layer2_outputs(6991);
    outputs(8052) <= layer2_outputs(7862);
    outputs(8053) <= not(layer2_outputs(4996));
    outputs(8054) <= not(layer2_outputs(5641));
    outputs(8055) <= layer2_outputs(9793);
    outputs(8056) <= layer2_outputs(5266);
    outputs(8057) <= not(layer2_outputs(3678)) or (layer2_outputs(826));
    outputs(8058) <= layer2_outputs(7961);
    outputs(8059) <= layer2_outputs(7649);
    outputs(8060) <= layer2_outputs(7885);
    outputs(8061) <= not((layer2_outputs(6626)) or (layer2_outputs(7650)));
    outputs(8062) <= not(layer2_outputs(1747));
    outputs(8063) <= not(layer2_outputs(9832));
    outputs(8064) <= not(layer2_outputs(9472));
    outputs(8065) <= layer2_outputs(2323);
    outputs(8066) <= not(layer2_outputs(4347));
    outputs(8067) <= (layer2_outputs(7456)) xor (layer2_outputs(7879));
    outputs(8068) <= not(layer2_outputs(7762));
    outputs(8069) <= (layer2_outputs(570)) and not (layer2_outputs(1654));
    outputs(8070) <= not(layer2_outputs(3404));
    outputs(8071) <= not(layer2_outputs(5963));
    outputs(8072) <= layer2_outputs(1561);
    outputs(8073) <= layer2_outputs(5748);
    outputs(8074) <= (layer2_outputs(5782)) and (layer2_outputs(7558));
    outputs(8075) <= layer2_outputs(768);
    outputs(8076) <= (layer2_outputs(1443)) xor (layer2_outputs(9850));
    outputs(8077) <= not((layer2_outputs(2476)) or (layer2_outputs(2167)));
    outputs(8078) <= not(layer2_outputs(4175));
    outputs(8079) <= (layer2_outputs(3432)) and (layer2_outputs(8795));
    outputs(8080) <= (layer2_outputs(5685)) xor (layer2_outputs(3524));
    outputs(8081) <= not(layer2_outputs(1774));
    outputs(8082) <= not((layer2_outputs(6564)) and (layer2_outputs(8938)));
    outputs(8083) <= layer2_outputs(2457);
    outputs(8084) <= not((layer2_outputs(6818)) xor (layer2_outputs(942)));
    outputs(8085) <= (layer2_outputs(4223)) xor (layer2_outputs(14));
    outputs(8086) <= layer2_outputs(1417);
    outputs(8087) <= layer2_outputs(7661);
    outputs(8088) <= not(layer2_outputs(1455));
    outputs(8089) <= layer2_outputs(3924);
    outputs(8090) <= not((layer2_outputs(3971)) or (layer2_outputs(4464)));
    outputs(8091) <= (layer2_outputs(1303)) and (layer2_outputs(7539));
    outputs(8092) <= layer2_outputs(7201);
    outputs(8093) <= not(layer2_outputs(7845));
    outputs(8094) <= not(layer2_outputs(9522));
    outputs(8095) <= not(layer2_outputs(6195));
    outputs(8096) <= not((layer2_outputs(985)) xor (layer2_outputs(3452)));
    outputs(8097) <= not(layer2_outputs(3125));
    outputs(8098) <= not(layer2_outputs(8343));
    outputs(8099) <= not((layer2_outputs(3664)) xor (layer2_outputs(3240)));
    outputs(8100) <= layer2_outputs(919);
    outputs(8101) <= layer2_outputs(1055);
    outputs(8102) <= layer2_outputs(4927);
    outputs(8103) <= layer2_outputs(5372);
    outputs(8104) <= not(layer2_outputs(10239)) or (layer2_outputs(7180));
    outputs(8105) <= not(layer2_outputs(9407));
    outputs(8106) <= layer2_outputs(4798);
    outputs(8107) <= layer2_outputs(6147);
    outputs(8108) <= not(layer2_outputs(1298));
    outputs(8109) <= not(layer2_outputs(1839));
    outputs(8110) <= layer2_outputs(121);
    outputs(8111) <= not(layer2_outputs(7370));
    outputs(8112) <= not(layer2_outputs(1965));
    outputs(8113) <= not((layer2_outputs(9391)) xor (layer2_outputs(5975)));
    outputs(8114) <= layer2_outputs(4322);
    outputs(8115) <= layer2_outputs(8058);
    outputs(8116) <= layer2_outputs(6128);
    outputs(8117) <= (layer2_outputs(5637)) or (layer2_outputs(2491));
    outputs(8118) <= layer2_outputs(3706);
    outputs(8119) <= (layer2_outputs(620)) xor (layer2_outputs(8183));
    outputs(8120) <= (layer2_outputs(7890)) and not (layer2_outputs(6137));
    outputs(8121) <= layer2_outputs(8164);
    outputs(8122) <= layer2_outputs(6510);
    outputs(8123) <= layer2_outputs(8268);
    outputs(8124) <= layer2_outputs(8303);
    outputs(8125) <= layer2_outputs(8963);
    outputs(8126) <= not((layer2_outputs(8093)) or (layer2_outputs(8625)));
    outputs(8127) <= not(layer2_outputs(4352));
    outputs(8128) <= layer2_outputs(6835);
    outputs(8129) <= layer2_outputs(4381);
    outputs(8130) <= layer2_outputs(6314);
    outputs(8131) <= (layer2_outputs(6681)) and not (layer2_outputs(8575));
    outputs(8132) <= layer2_outputs(1757);
    outputs(8133) <= not(layer2_outputs(6798));
    outputs(8134) <= not(layer2_outputs(6732));
    outputs(8135) <= not((layer2_outputs(9752)) xor (layer2_outputs(5922)));
    outputs(8136) <= not(layer2_outputs(2020));
    outputs(8137) <= layer2_outputs(8102);
    outputs(8138) <= layer2_outputs(8426);
    outputs(8139) <= (layer2_outputs(6611)) xor (layer2_outputs(4816));
    outputs(8140) <= not((layer2_outputs(6531)) xor (layer2_outputs(4737)));
    outputs(8141) <= (layer2_outputs(2187)) xor (layer2_outputs(6694));
    outputs(8142) <= not((layer2_outputs(1844)) or (layer2_outputs(3158)));
    outputs(8143) <= (layer2_outputs(4784)) xor (layer2_outputs(9165));
    outputs(8144) <= (layer2_outputs(708)) and (layer2_outputs(3919));
    outputs(8145) <= layer2_outputs(8359);
    outputs(8146) <= (layer2_outputs(4042)) xor (layer2_outputs(5099));
    outputs(8147) <= not(layer2_outputs(1037));
    outputs(8148) <= not(layer2_outputs(81));
    outputs(8149) <= not(layer2_outputs(3020));
    outputs(8150) <= layer2_outputs(4726);
    outputs(8151) <= not(layer2_outputs(1610));
    outputs(8152) <= (layer2_outputs(7553)) xor (layer2_outputs(2420));
    outputs(8153) <= not((layer2_outputs(8940)) and (layer2_outputs(7493)));
    outputs(8154) <= layer2_outputs(3185);
    outputs(8155) <= layer2_outputs(9175);
    outputs(8156) <= layer2_outputs(5018);
    outputs(8157) <= not(layer2_outputs(1812));
    outputs(8158) <= not(layer2_outputs(9104));
    outputs(8159) <= layer2_outputs(1491);
    outputs(8160) <= not((layer2_outputs(5415)) xor (layer2_outputs(6589)));
    outputs(8161) <= (layer2_outputs(6082)) xor (layer2_outputs(4282));
    outputs(8162) <= (layer2_outputs(6720)) and (layer2_outputs(8606));
    outputs(8163) <= (layer2_outputs(4739)) and (layer2_outputs(6817));
    outputs(8164) <= not(layer2_outputs(9871));
    outputs(8165) <= not((layer2_outputs(6994)) or (layer2_outputs(7513)));
    outputs(8166) <= not(layer2_outputs(5597));
    outputs(8167) <= not((layer2_outputs(6777)) xor (layer2_outputs(2224)));
    outputs(8168) <= (layer2_outputs(5509)) and (layer2_outputs(2922));
    outputs(8169) <= (layer2_outputs(9508)) and not (layer2_outputs(4878));
    outputs(8170) <= not(layer2_outputs(5566));
    outputs(8171) <= not(layer2_outputs(7926));
    outputs(8172) <= layer2_outputs(4556);
    outputs(8173) <= layer2_outputs(3896);
    outputs(8174) <= not(layer2_outputs(6630));
    outputs(8175) <= not((layer2_outputs(5603)) or (layer2_outputs(4251)));
    outputs(8176) <= not((layer2_outputs(6437)) xor (layer2_outputs(7799)));
    outputs(8177) <= layer2_outputs(2245);
    outputs(8178) <= (layer2_outputs(8763)) and not (layer2_outputs(9592));
    outputs(8179) <= not((layer2_outputs(3572)) xor (layer2_outputs(7153)));
    outputs(8180) <= not(layer2_outputs(1437));
    outputs(8181) <= not((layer2_outputs(1888)) or (layer2_outputs(7742)));
    outputs(8182) <= layer2_outputs(5846);
    outputs(8183) <= (layer2_outputs(3710)) and not (layer2_outputs(4873));
    outputs(8184) <= not(layer2_outputs(3537));
    outputs(8185) <= (layer2_outputs(1326)) xor (layer2_outputs(2582));
    outputs(8186) <= not((layer2_outputs(7828)) xor (layer2_outputs(6228)));
    outputs(8187) <= layer2_outputs(3942);
    outputs(8188) <= not(layer2_outputs(2022));
    outputs(8189) <= layer2_outputs(4322);
    outputs(8190) <= layer2_outputs(6116);
    outputs(8191) <= layer2_outputs(7977);
    outputs(8192) <= layer2_outputs(9061);
    outputs(8193) <= not((layer2_outputs(8704)) xor (layer2_outputs(3730)));
    outputs(8194) <= not((layer2_outputs(2600)) and (layer2_outputs(1960)));
    outputs(8195) <= not(layer2_outputs(3994));
    outputs(8196) <= not((layer2_outputs(4369)) xor (layer2_outputs(6732)));
    outputs(8197) <= layer2_outputs(3868);
    outputs(8198) <= not(layer2_outputs(1787)) or (layer2_outputs(9896));
    outputs(8199) <= not(layer2_outputs(5786)) or (layer2_outputs(9492));
    outputs(8200) <= not(layer2_outputs(5988)) or (layer2_outputs(7616));
    outputs(8201) <= (layer2_outputs(4211)) or (layer2_outputs(7530));
    outputs(8202) <= layer2_outputs(3758);
    outputs(8203) <= not((layer2_outputs(4149)) xor (layer2_outputs(9345)));
    outputs(8204) <= (layer2_outputs(3970)) and (layer2_outputs(9641));
    outputs(8205) <= not(layer2_outputs(1015));
    outputs(8206) <= (layer2_outputs(1630)) xor (layer2_outputs(4431));
    outputs(8207) <= not(layer2_outputs(5533));
    outputs(8208) <= layer2_outputs(5879);
    outputs(8209) <= not(layer2_outputs(925));
    outputs(8210) <= not((layer2_outputs(8167)) xor (layer2_outputs(9418)));
    outputs(8211) <= not((layer2_outputs(6467)) xor (layer2_outputs(9137)));
    outputs(8212) <= not(layer2_outputs(4637)) or (layer2_outputs(593));
    outputs(8213) <= not(layer2_outputs(1632)) or (layer2_outputs(5784));
    outputs(8214) <= not(layer2_outputs(389));
    outputs(8215) <= not(layer2_outputs(411)) or (layer2_outputs(4813));
    outputs(8216) <= not((layer2_outputs(7804)) xor (layer2_outputs(4680)));
    outputs(8217) <= not(layer2_outputs(7578));
    outputs(8218) <= layer2_outputs(3303);
    outputs(8219) <= not((layer2_outputs(9966)) xor (layer2_outputs(3730)));
    outputs(8220) <= not(layer2_outputs(6309));
    outputs(8221) <= not(layer2_outputs(4928));
    outputs(8222) <= layer2_outputs(4712);
    outputs(8223) <= layer2_outputs(2992);
    outputs(8224) <= layer2_outputs(4610);
    outputs(8225) <= (layer2_outputs(7134)) or (layer2_outputs(8612));
    outputs(8226) <= not(layer2_outputs(5611));
    outputs(8227) <= (layer2_outputs(1380)) xor (layer2_outputs(8789));
    outputs(8228) <= not((layer2_outputs(5089)) xor (layer2_outputs(6787)));
    outputs(8229) <= not(layer2_outputs(1383));
    outputs(8230) <= not((layer2_outputs(8828)) xor (layer2_outputs(5909)));
    outputs(8231) <= (layer2_outputs(8531)) or (layer2_outputs(4302));
    outputs(8232) <= layer2_outputs(9478);
    outputs(8233) <= layer2_outputs(7294);
    outputs(8234) <= (layer2_outputs(8479)) xor (layer2_outputs(5273));
    outputs(8235) <= not(layer2_outputs(6740));
    outputs(8236) <= not(layer2_outputs(4819)) or (layer2_outputs(1847));
    outputs(8237) <= not(layer2_outputs(489));
    outputs(8238) <= not((layer2_outputs(4475)) xor (layer2_outputs(8584)));
    outputs(8239) <= layer2_outputs(9597);
    outputs(8240) <= not(layer2_outputs(1398));
    outputs(8241) <= layer2_outputs(7312);
    outputs(8242) <= not(layer2_outputs(3553));
    outputs(8243) <= not(layer2_outputs(9960)) or (layer2_outputs(5248));
    outputs(8244) <= not(layer2_outputs(9105));
    outputs(8245) <= not(layer2_outputs(946));
    outputs(8246) <= not((layer2_outputs(5440)) xor (layer2_outputs(6970)));
    outputs(8247) <= layer2_outputs(2030);
    outputs(8248) <= not(layer2_outputs(2039));
    outputs(8249) <= (layer2_outputs(7231)) or (layer2_outputs(199));
    outputs(8250) <= not(layer2_outputs(8022));
    outputs(8251) <= not((layer2_outputs(3613)) xor (layer2_outputs(909)));
    outputs(8252) <= layer2_outputs(737);
    outputs(8253) <= layer2_outputs(3674);
    outputs(8254) <= not(layer2_outputs(7812)) or (layer2_outputs(9314));
    outputs(8255) <= (layer2_outputs(1809)) or (layer2_outputs(9223));
    outputs(8256) <= not(layer2_outputs(7315));
    outputs(8257) <= layer2_outputs(1130);
    outputs(8258) <= not(layer2_outputs(1905));
    outputs(8259) <= layer2_outputs(5262);
    outputs(8260) <= layer2_outputs(3518);
    outputs(8261) <= layer2_outputs(8072);
    outputs(8262) <= not((layer2_outputs(8279)) xor (layer2_outputs(7032)));
    outputs(8263) <= not((layer2_outputs(5389)) xor (layer2_outputs(7564)));
    outputs(8264) <= layer2_outputs(674);
    outputs(8265) <= (layer2_outputs(841)) xor (layer2_outputs(3883));
    outputs(8266) <= not(layer2_outputs(1240));
    outputs(8267) <= layer2_outputs(862);
    outputs(8268) <= (layer2_outputs(7489)) and not (layer2_outputs(5743));
    outputs(8269) <= layer2_outputs(6675);
    outputs(8270) <= not(layer2_outputs(9909));
    outputs(8271) <= not((layer2_outputs(8003)) xor (layer2_outputs(443)));
    outputs(8272) <= not((layer2_outputs(6773)) xor (layer2_outputs(7100)));
    outputs(8273) <= (layer2_outputs(5837)) xor (layer2_outputs(467));
    outputs(8274) <= (layer2_outputs(4159)) xor (layer2_outputs(7495));
    outputs(8275) <= not(layer2_outputs(1307));
    outputs(8276) <= layer2_outputs(147);
    outputs(8277) <= not((layer2_outputs(6037)) xor (layer2_outputs(1808)));
    outputs(8278) <= not((layer2_outputs(8961)) or (layer2_outputs(5665)));
    outputs(8279) <= (layer2_outputs(5324)) xor (layer2_outputs(6010));
    outputs(8280) <= not((layer2_outputs(6002)) or (layer2_outputs(8752)));
    outputs(8281) <= not(layer2_outputs(3115));
    outputs(8282) <= not(layer2_outputs(1729)) or (layer2_outputs(6070));
    outputs(8283) <= (layer2_outputs(10016)) xor (layer2_outputs(1657));
    outputs(8284) <= (layer2_outputs(875)) xor (layer2_outputs(6468));
    outputs(8285) <= not(layer2_outputs(4727));
    outputs(8286) <= (layer2_outputs(305)) and not (layer2_outputs(866));
    outputs(8287) <= (layer2_outputs(8748)) and (layer2_outputs(4960));
    outputs(8288) <= not((layer2_outputs(7582)) xor (layer2_outputs(6959)));
    outputs(8289) <= layer2_outputs(8642);
    outputs(8290) <= not(layer2_outputs(8179));
    outputs(8291) <= not(layer2_outputs(2594)) or (layer2_outputs(167));
    outputs(8292) <= not(layer2_outputs(3874));
    outputs(8293) <= (layer2_outputs(740)) xor (layer2_outputs(5087));
    outputs(8294) <= not((layer2_outputs(391)) xor (layer2_outputs(9638)));
    outputs(8295) <= '1';
    outputs(8296) <= not(layer2_outputs(2779));
    outputs(8297) <= layer2_outputs(2524);
    outputs(8298) <= (layer2_outputs(5754)) xor (layer2_outputs(6569));
    outputs(8299) <= (layer2_outputs(1357)) xor (layer2_outputs(9857));
    outputs(8300) <= (layer2_outputs(75)) xor (layer2_outputs(1773));
    outputs(8301) <= not((layer2_outputs(1713)) and (layer2_outputs(2984)));
    outputs(8302) <= layer2_outputs(8261);
    outputs(8303) <= (layer2_outputs(2418)) xor (layer2_outputs(2291));
    outputs(8304) <= layer2_outputs(5163);
    outputs(8305) <= (layer2_outputs(10076)) or (layer2_outputs(1812));
    outputs(8306) <= not((layer2_outputs(3222)) xor (layer2_outputs(9398)));
    outputs(8307) <= (layer2_outputs(6502)) xor (layer2_outputs(6531));
    outputs(8308) <= layer2_outputs(8893);
    outputs(8309) <= not(layer2_outputs(1453));
    outputs(8310) <= not((layer2_outputs(7735)) or (layer2_outputs(2696)));
    outputs(8311) <= (layer2_outputs(8523)) xor (layer2_outputs(9028));
    outputs(8312) <= (layer2_outputs(1013)) xor (layer2_outputs(1568));
    outputs(8313) <= not(layer2_outputs(6721));
    outputs(8314) <= (layer2_outputs(9099)) xor (layer2_outputs(3150));
    outputs(8315) <= (layer2_outputs(8815)) xor (layer2_outputs(7408));
    outputs(8316) <= not(layer2_outputs(9336));
    outputs(8317) <= layer2_outputs(4519);
    outputs(8318) <= layer2_outputs(6884);
    outputs(8319) <= (layer2_outputs(3660)) xor (layer2_outputs(652));
    outputs(8320) <= not(layer2_outputs(9069)) or (layer2_outputs(8550));
    outputs(8321) <= (layer2_outputs(6247)) and not (layer2_outputs(9646));
    outputs(8322) <= not(layer2_outputs(4275));
    outputs(8323) <= not((layer2_outputs(9712)) xor (layer2_outputs(7027)));
    outputs(8324) <= not((layer2_outputs(9448)) and (layer2_outputs(2733)));
    outputs(8325) <= not(layer2_outputs(1186));
    outputs(8326) <= layer2_outputs(9067);
    outputs(8327) <= not(layer2_outputs(3802)) or (layer2_outputs(8503));
    outputs(8328) <= not((layer2_outputs(7232)) xor (layer2_outputs(9)));
    outputs(8329) <= not((layer2_outputs(1780)) and (layer2_outputs(7933)));
    outputs(8330) <= (layer2_outputs(8634)) and not (layer2_outputs(6298));
    outputs(8331) <= (layer2_outputs(3164)) xor (layer2_outputs(3145));
    outputs(8332) <= (layer2_outputs(6536)) xor (layer2_outputs(1234));
    outputs(8333) <= (layer2_outputs(5177)) xor (layer2_outputs(2297));
    outputs(8334) <= not(layer2_outputs(3369));
    outputs(8335) <= not(layer2_outputs(3111)) or (layer2_outputs(1884));
    outputs(8336) <= layer2_outputs(1711);
    outputs(8337) <= not((layer2_outputs(2308)) xor (layer2_outputs(5845)));
    outputs(8338) <= (layer2_outputs(4203)) and (layer2_outputs(3707));
    outputs(8339) <= not(layer2_outputs(9738));
    outputs(8340) <= layer2_outputs(1297);
    outputs(8341) <= not(layer2_outputs(10235)) or (layer2_outputs(6858));
    outputs(8342) <= not((layer2_outputs(436)) xor (layer2_outputs(1793)));
    outputs(8343) <= not(layer2_outputs(4828));
    outputs(8344) <= not(layer2_outputs(3965)) or (layer2_outputs(179));
    outputs(8345) <= layer2_outputs(8791);
    outputs(8346) <= (layer2_outputs(4671)) or (layer2_outputs(9075));
    outputs(8347) <= not(layer2_outputs(6807));
    outputs(8348) <= not(layer2_outputs(9728));
    outputs(8349) <= (layer2_outputs(6776)) xor (layer2_outputs(8786));
    outputs(8350) <= not(layer2_outputs(9921)) or (layer2_outputs(8620));
    outputs(8351) <= layer2_outputs(1728);
    outputs(8352) <= (layer2_outputs(4287)) xor (layer2_outputs(9143));
    outputs(8353) <= layer2_outputs(2139);
    outputs(8354) <= layer2_outputs(355);
    outputs(8355) <= (layer2_outputs(7963)) and not (layer2_outputs(3100));
    outputs(8356) <= layer2_outputs(874);
    outputs(8357) <= not(layer2_outputs(2279));
    outputs(8358) <= (layer2_outputs(2529)) xor (layer2_outputs(7117));
    outputs(8359) <= (layer2_outputs(5204)) xor (layer2_outputs(7216));
    outputs(8360) <= layer2_outputs(2791);
    outputs(8361) <= (layer2_outputs(1933)) xor (layer2_outputs(3975));
    outputs(8362) <= not(layer2_outputs(7145));
    outputs(8363) <= layer2_outputs(7042);
    outputs(8364) <= layer2_outputs(4413);
    outputs(8365) <= (layer2_outputs(4610)) and not (layer2_outputs(2258));
    outputs(8366) <= (layer2_outputs(4543)) xor (layer2_outputs(2340));
    outputs(8367) <= not(layer2_outputs(8468));
    outputs(8368) <= not(layer2_outputs(9940));
    outputs(8369) <= layer2_outputs(2461);
    outputs(8370) <= not(layer2_outputs(8112));
    outputs(8371) <= layer2_outputs(2335);
    outputs(8372) <= not(layer2_outputs(5621));
    outputs(8373) <= (layer2_outputs(5716)) and not (layer2_outputs(1523));
    outputs(8374) <= (layer2_outputs(1489)) or (layer2_outputs(9011));
    outputs(8375) <= not(layer2_outputs(6717));
    outputs(8376) <= layer2_outputs(554);
    outputs(8377) <= not(layer2_outputs(1036));
    outputs(8378) <= not(layer2_outputs(1632)) or (layer2_outputs(5411));
    outputs(8379) <= not((layer2_outputs(8970)) xor (layer2_outputs(8240)));
    outputs(8380) <= not((layer2_outputs(4592)) and (layer2_outputs(5088)));
    outputs(8381) <= layer2_outputs(2765);
    outputs(8382) <= not((layer2_outputs(735)) xor (layer2_outputs(9199)));
    outputs(8383) <= layer2_outputs(1000);
    outputs(8384) <= layer2_outputs(2572);
    outputs(8385) <= not(layer2_outputs(8905));
    outputs(8386) <= (layer2_outputs(3644)) and not (layer2_outputs(691));
    outputs(8387) <= not(layer2_outputs(2272));
    outputs(8388) <= layer2_outputs(2485);
    outputs(8389) <= not(layer2_outputs(5007));
    outputs(8390) <= not(layer2_outputs(4951));
    outputs(8391) <= not(layer2_outputs(104));
    outputs(8392) <= (layer2_outputs(2310)) or (layer2_outputs(8502));
    outputs(8393) <= (layer2_outputs(2674)) xor (layer2_outputs(635));
    outputs(8394) <= layer2_outputs(2658);
    outputs(8395) <= (layer2_outputs(2141)) xor (layer2_outputs(205));
    outputs(8396) <= (layer2_outputs(513)) or (layer2_outputs(1733));
    outputs(8397) <= layer2_outputs(1824);
    outputs(8398) <= (layer2_outputs(105)) xor (layer2_outputs(10067));
    outputs(8399) <= not(layer2_outputs(5647));
    outputs(8400) <= not((layer2_outputs(4377)) xor (layer2_outputs(4017)));
    outputs(8401) <= not((layer2_outputs(4752)) xor (layer2_outputs(7240)));
    outputs(8402) <= (layer2_outputs(1567)) xor (layer2_outputs(7746));
    outputs(8403) <= not(layer2_outputs(5440)) or (layer2_outputs(3221));
    outputs(8404) <= layer2_outputs(8979);
    outputs(8405) <= (layer2_outputs(9217)) or (layer2_outputs(9461));
    outputs(8406) <= not((layer2_outputs(2284)) or (layer2_outputs(7956)));
    outputs(8407) <= not((layer2_outputs(7513)) xor (layer2_outputs(1322)));
    outputs(8408) <= not((layer2_outputs(7958)) xor (layer2_outputs(8706)));
    outputs(8409) <= not((layer2_outputs(111)) xor (layer2_outputs(1569)));
    outputs(8410) <= not(layer2_outputs(3750));
    outputs(8411) <= (layer2_outputs(193)) xor (layer2_outputs(3609));
    outputs(8412) <= (layer2_outputs(1519)) xor (layer2_outputs(8734));
    outputs(8413) <= not((layer2_outputs(7638)) xor (layer2_outputs(2718)));
    outputs(8414) <= not(layer2_outputs(5235));
    outputs(8415) <= not(layer2_outputs(9233)) or (layer2_outputs(9159));
    outputs(8416) <= not(layer2_outputs(2533)) or (layer2_outputs(5163));
    outputs(8417) <= (layer2_outputs(681)) xor (layer2_outputs(9890));
    outputs(8418) <= layer2_outputs(3026);
    outputs(8419) <= not(layer2_outputs(3269));
    outputs(8420) <= not((layer2_outputs(2978)) xor (layer2_outputs(1624)));
    outputs(8421) <= not((layer2_outputs(5506)) xor (layer2_outputs(5675)));
    outputs(8422) <= (layer2_outputs(5346)) xor (layer2_outputs(1762));
    outputs(8423) <= layer2_outputs(4038);
    outputs(8424) <= (layer2_outputs(1753)) xor (layer2_outputs(7683));
    outputs(8425) <= (layer2_outputs(1926)) or (layer2_outputs(4374));
    outputs(8426) <= not((layer2_outputs(4035)) xor (layer2_outputs(9699)));
    outputs(8427) <= layer2_outputs(658);
    outputs(8428) <= (layer2_outputs(2429)) xor (layer2_outputs(1893));
    outputs(8429) <= not((layer2_outputs(2423)) and (layer2_outputs(621)));
    outputs(8430) <= not((layer2_outputs(9906)) or (layer2_outputs(2612)));
    outputs(8431) <= not(layer2_outputs(4419));
    outputs(8432) <= layer2_outputs(3653);
    outputs(8433) <= (layer2_outputs(7026)) xor (layer2_outputs(1280));
    outputs(8434) <= not(layer2_outputs(7351));
    outputs(8435) <= layer2_outputs(3992);
    outputs(8436) <= layer2_outputs(4292);
    outputs(8437) <= not((layer2_outputs(7832)) xor (layer2_outputs(7907)));
    outputs(8438) <= not(layer2_outputs(5323));
    outputs(8439) <= layer2_outputs(3542);
    outputs(8440) <= not((layer2_outputs(8433)) xor (layer2_outputs(8715)));
    outputs(8441) <= not(layer2_outputs(9887));
    outputs(8442) <= (layer2_outputs(2994)) xor (layer2_outputs(2938));
    outputs(8443) <= layer2_outputs(319);
    outputs(8444) <= not(layer2_outputs(5652)) or (layer2_outputs(6383));
    outputs(8445) <= not(layer2_outputs(8992));
    outputs(8446) <= not(layer2_outputs(4428));
    outputs(8447) <= (layer2_outputs(3595)) xor (layer2_outputs(4446));
    outputs(8448) <= layer2_outputs(6516);
    outputs(8449) <= not((layer2_outputs(2953)) xor (layer2_outputs(9733)));
    outputs(8450) <= not(layer2_outputs(5139));
    outputs(8451) <= not((layer2_outputs(9813)) xor (layer2_outputs(7548)));
    outputs(8452) <= (layer2_outputs(6717)) xor (layer2_outputs(3677));
    outputs(8453) <= not((layer2_outputs(6966)) or (layer2_outputs(7003)));
    outputs(8454) <= not(layer2_outputs(8182));
    outputs(8455) <= (layer2_outputs(9251)) and not (layer2_outputs(6025));
    outputs(8456) <= not(layer2_outputs(9088)) or (layer2_outputs(4729));
    outputs(8457) <= not((layer2_outputs(8907)) xor (layer2_outputs(8074)));
    outputs(8458) <= layer2_outputs(450);
    outputs(8459) <= not((layer2_outputs(9659)) and (layer2_outputs(8399)));
    outputs(8460) <= (layer2_outputs(1300)) or (layer2_outputs(9871));
    outputs(8461) <= (layer2_outputs(5683)) xor (layer2_outputs(6573));
    outputs(8462) <= layer2_outputs(2480);
    outputs(8463) <= (layer2_outputs(2236)) xor (layer2_outputs(2041));
    outputs(8464) <= not((layer2_outputs(4277)) xor (layer2_outputs(3327)));
    outputs(8465) <= not((layer2_outputs(2285)) xor (layer2_outputs(7259)));
    outputs(8466) <= not((layer2_outputs(8855)) and (layer2_outputs(787)));
    outputs(8467) <= layer2_outputs(1524);
    outputs(8468) <= (layer2_outputs(8762)) or (layer2_outputs(2845));
    outputs(8469) <= (layer2_outputs(9785)) or (layer2_outputs(10189));
    outputs(8470) <= not((layer2_outputs(1093)) xor (layer2_outputs(3555)));
    outputs(8471) <= not(layer2_outputs(8805));
    outputs(8472) <= (layer2_outputs(3600)) xor (layer2_outputs(9802));
    outputs(8473) <= (layer2_outputs(556)) and not (layer2_outputs(741));
    outputs(8474) <= not((layer2_outputs(7948)) and (layer2_outputs(869)));
    outputs(8475) <= not((layer2_outputs(5651)) xor (layer2_outputs(6824)));
    outputs(8476) <= not(layer2_outputs(58));
    outputs(8477) <= not((layer2_outputs(9101)) xor (layer2_outputs(7095)));
    outputs(8478) <= layer2_outputs(10158);
    outputs(8479) <= layer2_outputs(1716);
    outputs(8480) <= (layer2_outputs(4181)) xor (layer2_outputs(2408));
    outputs(8481) <= (layer2_outputs(3708)) and not (layer2_outputs(3543));
    outputs(8482) <= (layer2_outputs(3211)) xor (layer2_outputs(4115));
    outputs(8483) <= (layer2_outputs(9689)) xor (layer2_outputs(840));
    outputs(8484) <= not(layer2_outputs(9562));
    outputs(8485) <= not(layer2_outputs(4536));
    outputs(8486) <= not(layer2_outputs(1475));
    outputs(8487) <= not(layer2_outputs(1047));
    outputs(8488) <= not(layer2_outputs(6042));
    outputs(8489) <= not(layer2_outputs(5172)) or (layer2_outputs(6776));
    outputs(8490) <= layer2_outputs(233);
    outputs(8491) <= not(layer2_outputs(9797)) or (layer2_outputs(6455));
    outputs(8492) <= not((layer2_outputs(2313)) xor (layer2_outputs(5103)));
    outputs(8493) <= (layer2_outputs(1041)) xor (layer2_outputs(4099));
    outputs(8494) <= layer2_outputs(7954);
    outputs(8495) <= layer2_outputs(7917);
    outputs(8496) <= not(layer2_outputs(4537)) or (layer2_outputs(6573));
    outputs(8497) <= (layer2_outputs(4712)) and not (layer2_outputs(3563));
    outputs(8498) <= not(layer2_outputs(1569));
    outputs(8499) <= (layer2_outputs(9191)) xor (layer2_outputs(656));
    outputs(8500) <= not(layer2_outputs(3315)) or (layer2_outputs(8193));
    outputs(8501) <= layer2_outputs(967);
    outputs(8502) <= (layer2_outputs(1309)) xor (layer2_outputs(220));
    outputs(8503) <= layer2_outputs(1447);
    outputs(8504) <= (layer2_outputs(6925)) xor (layer2_outputs(6180));
    outputs(8505) <= not((layer2_outputs(2090)) xor (layer2_outputs(4243)));
    outputs(8506) <= (layer2_outputs(7878)) xor (layer2_outputs(6638));
    outputs(8507) <= not((layer2_outputs(9721)) xor (layer2_outputs(5970)));
    outputs(8508) <= (layer2_outputs(8)) xor (layer2_outputs(2749));
    outputs(8509) <= not(layer2_outputs(85)) or (layer2_outputs(4027));
    outputs(8510) <= not((layer2_outputs(9117)) xor (layer2_outputs(7454)));
    outputs(8511) <= not((layer2_outputs(8740)) xor (layer2_outputs(4844)));
    outputs(8512) <= layer2_outputs(5694);
    outputs(8513) <= not((layer2_outputs(3648)) and (layer2_outputs(7313)));
    outputs(8514) <= not(layer2_outputs(934));
    outputs(8515) <= (layer2_outputs(6129)) xor (layer2_outputs(5514));
    outputs(8516) <= layer2_outputs(5366);
    outputs(8517) <= (layer2_outputs(9121)) xor (layer2_outputs(10026));
    outputs(8518) <= layer2_outputs(1871);
    outputs(8519) <= layer2_outputs(10188);
    outputs(8520) <= layer2_outputs(9845);
    outputs(8521) <= not(layer2_outputs(9827));
    outputs(8522) <= not(layer2_outputs(6868)) or (layer2_outputs(2852));
    outputs(8523) <= not(layer2_outputs(5589));
    outputs(8524) <= not(layer2_outputs(9950)) or (layer2_outputs(10026));
    outputs(8525) <= not((layer2_outputs(8389)) xor (layer2_outputs(4438)));
    outputs(8526) <= not((layer2_outputs(8042)) xor (layer2_outputs(2417)));
    outputs(8527) <= (layer2_outputs(2874)) xor (layer2_outputs(8830));
    outputs(8528) <= (layer2_outputs(5277)) xor (layer2_outputs(1672));
    outputs(8529) <= not(layer2_outputs(8969));
    outputs(8530) <= layer2_outputs(4718);
    outputs(8531) <= (layer2_outputs(2302)) xor (layer2_outputs(7441));
    outputs(8532) <= not(layer2_outputs(5583));
    outputs(8533) <= not((layer2_outputs(3522)) and (layer2_outputs(127)));
    outputs(8534) <= (layer2_outputs(8250)) xor (layer2_outputs(3030));
    outputs(8535) <= layer2_outputs(5820);
    outputs(8536) <= not(layer2_outputs(7676));
    outputs(8537) <= not(layer2_outputs(8733));
    outputs(8538) <= not((layer2_outputs(3852)) xor (layer2_outputs(5122)));
    outputs(8539) <= layer2_outputs(124);
    outputs(8540) <= layer2_outputs(10156);
    outputs(8541) <= not((layer2_outputs(7487)) and (layer2_outputs(5248)));
    outputs(8542) <= not((layer2_outputs(9747)) xor (layer2_outputs(2988)));
    outputs(8543) <= not(layer2_outputs(3512));
    outputs(8544) <= not(layer2_outputs(825));
    outputs(8545) <= not(layer2_outputs(8701));
    outputs(8546) <= not(layer2_outputs(6836)) or (layer2_outputs(2482));
    outputs(8547) <= layer2_outputs(743);
    outputs(8548) <= not((layer2_outputs(4909)) xor (layer2_outputs(4396)));
    outputs(8549) <= layer2_outputs(6919);
    outputs(8550) <= not((layer2_outputs(1992)) xor (layer2_outputs(4696)));
    outputs(8551) <= not((layer2_outputs(3463)) xor (layer2_outputs(9361)));
    outputs(8552) <= not(layer2_outputs(3885));
    outputs(8553) <= not(layer2_outputs(5960));
    outputs(8554) <= not((layer2_outputs(4583)) and (layer2_outputs(3227)));
    outputs(8555) <= (layer2_outputs(7780)) xor (layer2_outputs(8933));
    outputs(8556) <= layer2_outputs(1138);
    outputs(8557) <= not((layer2_outputs(969)) and (layer2_outputs(609)));
    outputs(8558) <= not(layer2_outputs(1978));
    outputs(8559) <= not(layer2_outputs(7555));
    outputs(8560) <= layer2_outputs(1891);
    outputs(8561) <= layer2_outputs(2460);
    outputs(8562) <= not(layer2_outputs(4831)) or (layer2_outputs(6295));
    outputs(8563) <= not(layer2_outputs(2787)) or (layer2_outputs(4972));
    outputs(8564) <= layer2_outputs(2117);
    outputs(8565) <= not((layer2_outputs(2681)) and (layer2_outputs(9985)));
    outputs(8566) <= not(layer2_outputs(8671));
    outputs(8567) <= not(layer2_outputs(7937));
    outputs(8568) <= (layer2_outputs(6680)) xor (layer2_outputs(9155));
    outputs(8569) <= (layer2_outputs(8346)) and not (layer2_outputs(5230));
    outputs(8570) <= layer2_outputs(4178);
    outputs(8571) <= layer2_outputs(1594);
    outputs(8572) <= layer2_outputs(8968);
    outputs(8573) <= (layer2_outputs(4669)) xor (layer2_outputs(6598));
    outputs(8574) <= (layer2_outputs(7132)) xor (layer2_outputs(3552));
    outputs(8575) <= not(layer2_outputs(8450));
    outputs(8576) <= not((layer2_outputs(7906)) xor (layer2_outputs(1294)));
    outputs(8577) <= not(layer2_outputs(5491));
    outputs(8578) <= layer2_outputs(4347);
    outputs(8579) <= not(layer2_outputs(3359)) or (layer2_outputs(920));
    outputs(8580) <= layer2_outputs(1623);
    outputs(8581) <= layer2_outputs(2068);
    outputs(8582) <= not((layer2_outputs(6484)) xor (layer2_outputs(5304)));
    outputs(8583) <= (layer2_outputs(5457)) and not (layer2_outputs(3322));
    outputs(8584) <= not(layer2_outputs(916));
    outputs(8585) <= not(layer2_outputs(3273));
    outputs(8586) <= not(layer2_outputs(7597));
    outputs(8587) <= layer2_outputs(5806);
    outputs(8588) <= layer2_outputs(214);
    outputs(8589) <= not((layer2_outputs(7168)) or (layer2_outputs(3416)));
    outputs(8590) <= layer2_outputs(7187);
    outputs(8591) <= (layer2_outputs(5336)) xor (layer2_outputs(899));
    outputs(8592) <= not(layer2_outputs(8405)) or (layer2_outputs(2415));
    outputs(8593) <= not(layer2_outputs(5127)) or (layer2_outputs(9786));
    outputs(8594) <= not(layer2_outputs(3385));
    outputs(8595) <= not((layer2_outputs(4505)) xor (layer2_outputs(2287)));
    outputs(8596) <= layer2_outputs(49);
    outputs(8597) <= layer2_outputs(4028);
    outputs(8598) <= not((layer2_outputs(8933)) xor (layer2_outputs(4667)));
    outputs(8599) <= (layer2_outputs(6556)) and not (layer2_outputs(977));
    outputs(8600) <= not(layer2_outputs(303));
    outputs(8601) <= layer2_outputs(1818);
    outputs(8602) <= (layer2_outputs(7189)) xor (layer2_outputs(4066));
    outputs(8603) <= not(layer2_outputs(838));
    outputs(8604) <= not(layer2_outputs(1878)) or (layer2_outputs(6585));
    outputs(8605) <= '1';
    outputs(8606) <= not(layer2_outputs(7685)) or (layer2_outputs(8478));
    outputs(8607) <= layer2_outputs(3956);
    outputs(8608) <= (layer2_outputs(1265)) xor (layer2_outputs(7844));
    outputs(8609) <= not(layer2_outputs(6182));
    outputs(8610) <= layer2_outputs(6441);
    outputs(8611) <= (layer2_outputs(3054)) and not (layer2_outputs(7586));
    outputs(8612) <= not((layer2_outputs(5012)) xor (layer2_outputs(143)));
    outputs(8613) <= layer2_outputs(6662);
    outputs(8614) <= layer2_outputs(314);
    outputs(8615) <= not(layer2_outputs(2286));
    outputs(8616) <= layer2_outputs(6871);
    outputs(8617) <= (layer2_outputs(8089)) and not (layer2_outputs(4332));
    outputs(8618) <= not((layer2_outputs(2133)) xor (layer2_outputs(5212)));
    outputs(8619) <= (layer2_outputs(8893)) xor (layer2_outputs(1505));
    outputs(8620) <= layer2_outputs(2667);
    outputs(8621) <= not(layer2_outputs(151));
    outputs(8622) <= not(layer2_outputs(5108));
    outputs(8623) <= (layer2_outputs(6709)) xor (layer2_outputs(5320));
    outputs(8624) <= layer2_outputs(3944);
    outputs(8625) <= (layer2_outputs(6491)) xor (layer2_outputs(7854));
    outputs(8626) <= not(layer2_outputs(2893));
    outputs(8627) <= (layer2_outputs(6323)) xor (layer2_outputs(3182));
    outputs(8628) <= not((layer2_outputs(637)) and (layer2_outputs(5302)));
    outputs(8629) <= not((layer2_outputs(6635)) and (layer2_outputs(4936)));
    outputs(8630) <= not((layer2_outputs(334)) xor (layer2_outputs(7991)));
    outputs(8631) <= (layer2_outputs(2535)) xor (layer2_outputs(9829));
    outputs(8632) <= (layer2_outputs(8097)) xor (layer2_outputs(803));
    outputs(8633) <= (layer2_outputs(3826)) xor (layer2_outputs(7157));
    outputs(8634) <= not(layer2_outputs(9903));
    outputs(8635) <= (layer2_outputs(9504)) and not (layer2_outputs(1918));
    outputs(8636) <= not(layer2_outputs(462));
    outputs(8637) <= layer2_outputs(1096);
    outputs(8638) <= layer2_outputs(3520);
    outputs(8639) <= layer2_outputs(6718);
    outputs(8640) <= not((layer2_outputs(9466)) xor (layer2_outputs(508)));
    outputs(8641) <= layer2_outputs(3752);
    outputs(8642) <= not(layer2_outputs(2664));
    outputs(8643) <= layer2_outputs(9184);
    outputs(8644) <= not((layer2_outputs(9392)) xor (layer2_outputs(9177)));
    outputs(8645) <= (layer2_outputs(5890)) xor (layer2_outputs(6394));
    outputs(8646) <= (layer2_outputs(2065)) xor (layer2_outputs(10057));
    outputs(8647) <= not(layer2_outputs(8035));
    outputs(8648) <= (layer2_outputs(1805)) xor (layer2_outputs(6476));
    outputs(8649) <= not((layer2_outputs(7299)) and (layer2_outputs(3957)));
    outputs(8650) <= not(layer2_outputs(2514));
    outputs(8651) <= (layer2_outputs(2948)) and not (layer2_outputs(3823));
    outputs(8652) <= not(layer2_outputs(8318));
    outputs(8653) <= layer2_outputs(2587);
    outputs(8654) <= not(layer2_outputs(8492));
    outputs(8655) <= not((layer2_outputs(2033)) xor (layer2_outputs(8421)));
    outputs(8656) <= layer2_outputs(5999);
    outputs(8657) <= (layer2_outputs(4825)) and not (layer2_outputs(4426));
    outputs(8658) <= (layer2_outputs(2742)) xor (layer2_outputs(1760));
    outputs(8659) <= not(layer2_outputs(8682));
    outputs(8660) <= (layer2_outputs(5464)) xor (layer2_outputs(1258));
    outputs(8661) <= not(layer2_outputs(5284));
    outputs(8662) <= not(layer2_outputs(10165)) or (layer2_outputs(2778));
    outputs(8663) <= not(layer2_outputs(7152));
    outputs(8664) <= (layer2_outputs(284)) xor (layer2_outputs(2571));
    outputs(8665) <= (layer2_outputs(7765)) xor (layer2_outputs(6591));
    outputs(8666) <= layer2_outputs(1466);
    outputs(8667) <= layer2_outputs(2882);
    outputs(8668) <= not((layer2_outputs(3285)) and (layer2_outputs(8219)));
    outputs(8669) <= layer2_outputs(4851);
    outputs(8670) <= not((layer2_outputs(1174)) xor (layer2_outputs(2237)));
    outputs(8671) <= not(layer2_outputs(7113));
    outputs(8672) <= not((layer2_outputs(5491)) xor (layer2_outputs(1150)));
    outputs(8673) <= not(layer2_outputs(3157));
    outputs(8674) <= layer2_outputs(9084);
    outputs(8675) <= (layer2_outputs(8887)) xor (layer2_outputs(6500));
    outputs(8676) <= not(layer2_outputs(3964));
    outputs(8677) <= layer2_outputs(7476);
    outputs(8678) <= not(layer2_outputs(1100));
    outputs(8679) <= not(layer2_outputs(3059)) or (layer2_outputs(3997));
    outputs(8680) <= (layer2_outputs(2593)) xor (layer2_outputs(8314));
    outputs(8681) <= not(layer2_outputs(1496));
    outputs(8682) <= not((layer2_outputs(3651)) xor (layer2_outputs(6811)));
    outputs(8683) <= not((layer2_outputs(6996)) xor (layer2_outputs(4468)));
    outputs(8684) <= not((layer2_outputs(921)) xor (layer2_outputs(6554)));
    outputs(8685) <= not(layer2_outputs(5448)) or (layer2_outputs(1903));
    outputs(8686) <= not(layer2_outputs(1576)) or (layer2_outputs(22));
    outputs(8687) <= not(layer2_outputs(7690));
    outputs(8688) <= layer2_outputs(7024);
    outputs(8689) <= not(layer2_outputs(2864));
    outputs(8690) <= not((layer2_outputs(2376)) and (layer2_outputs(9100)));
    outputs(8691) <= not(layer2_outputs(7874));
    outputs(8692) <= not((layer2_outputs(6177)) xor (layer2_outputs(1097)));
    outputs(8693) <= (layer2_outputs(3449)) xor (layer2_outputs(6710));
    outputs(8694) <= not((layer2_outputs(4333)) xor (layer2_outputs(4259)));
    outputs(8695) <= not((layer2_outputs(4521)) xor (layer2_outputs(8257)));
    outputs(8696) <= not(layer2_outputs(8607));
    outputs(8697) <= layer2_outputs(7327);
    outputs(8698) <= not(layer2_outputs(936));
    outputs(8699) <= not(layer2_outputs(8708)) or (layer2_outputs(7630));
    outputs(8700) <= layer2_outputs(86);
    outputs(8701) <= not(layer2_outputs(1650));
    outputs(8702) <= not(layer2_outputs(9310));
    outputs(8703) <= not(layer2_outputs(5923));
    outputs(8704) <= not(layer2_outputs(2031));
    outputs(8705) <= (layer2_outputs(293)) or (layer2_outputs(8288));
    outputs(8706) <= layer2_outputs(8860);
    outputs(8707) <= not((layer2_outputs(7401)) xor (layer2_outputs(9925)));
    outputs(8708) <= not((layer2_outputs(9194)) xor (layer2_outputs(7162)));
    outputs(8709) <= not(layer2_outputs(9150)) or (layer2_outputs(4340));
    outputs(8710) <= not(layer2_outputs(3705)) or (layer2_outputs(8881));
    outputs(8711) <= not((layer2_outputs(7982)) xor (layer2_outputs(6654)));
    outputs(8712) <= (layer2_outputs(5495)) xor (layer2_outputs(7193));
    outputs(8713) <= not(layer2_outputs(5745));
    outputs(8714) <= layer2_outputs(5283);
    outputs(8715) <= (layer2_outputs(6051)) xor (layer2_outputs(1005));
    outputs(8716) <= not(layer2_outputs(6661));
    outputs(8717) <= not((layer2_outputs(8745)) xor (layer2_outputs(3511)));
    outputs(8718) <= not(layer2_outputs(5220));
    outputs(8719) <= not(layer2_outputs(6165)) or (layer2_outputs(10008));
    outputs(8720) <= layer2_outputs(1772);
    outputs(8721) <= not((layer2_outputs(1325)) xor (layer2_outputs(994)));
    outputs(8722) <= not(layer2_outputs(8266));
    outputs(8723) <= layer2_outputs(134);
    outputs(8724) <= (layer2_outputs(2521)) and (layer2_outputs(7077));
    outputs(8725) <= not(layer2_outputs(989)) or (layer2_outputs(2731));
    outputs(8726) <= (layer2_outputs(8072)) xor (layer2_outputs(1242));
    outputs(8727) <= not(layer2_outputs(5803));
    outputs(8728) <= layer2_outputs(4721);
    outputs(8729) <= layer2_outputs(8478);
    outputs(8730) <= not(layer2_outputs(1694)) or (layer2_outputs(8982));
    outputs(8731) <= not((layer2_outputs(1622)) xor (layer2_outputs(357)));
    outputs(8732) <= not((layer2_outputs(1172)) and (layer2_outputs(391)));
    outputs(8733) <= layer2_outputs(3297);
    outputs(8734) <= not(layer2_outputs(6420));
    outputs(8735) <= layer2_outputs(6471);
    outputs(8736) <= not(layer2_outputs(1470));
    outputs(8737) <= (layer2_outputs(1088)) xor (layer2_outputs(9188));
    outputs(8738) <= layer2_outputs(7710);
    outputs(8739) <= not((layer2_outputs(7677)) or (layer2_outputs(2358)));
    outputs(8740) <= not(layer2_outputs(5263));
    outputs(8741) <= layer2_outputs(534);
    outputs(8742) <= not(layer2_outputs(6663));
    outputs(8743) <= not((layer2_outputs(4799)) and (layer2_outputs(1080)));
    outputs(8744) <= not((layer2_outputs(6903)) xor (layer2_outputs(2111)));
    outputs(8745) <= not((layer2_outputs(10183)) and (layer2_outputs(3522)));
    outputs(8746) <= layer2_outputs(6440);
    outputs(8747) <= not((layer2_outputs(6542)) xor (layer2_outputs(6041)));
    outputs(8748) <= layer2_outputs(8023);
    outputs(8749) <= not((layer2_outputs(4386)) xor (layer2_outputs(3112)));
    outputs(8750) <= (layer2_outputs(9485)) and (layer2_outputs(6039));
    outputs(8751) <= (layer2_outputs(4085)) xor (layer2_outputs(7257));
    outputs(8752) <= not((layer2_outputs(3830)) and (layer2_outputs(8633)));
    outputs(8753) <= layer2_outputs(10087);
    outputs(8754) <= (layer2_outputs(8514)) and not (layer2_outputs(7654));
    outputs(8755) <= layer2_outputs(9064);
    outputs(8756) <= (layer2_outputs(3722)) and not (layer2_outputs(2719));
    outputs(8757) <= layer2_outputs(8323);
    outputs(8758) <= not(layer2_outputs(2398)) or (layer2_outputs(9184));
    outputs(8759) <= (layer2_outputs(1675)) xor (layer2_outputs(5591));
    outputs(8760) <= layer2_outputs(7990);
    outputs(8761) <= not(layer2_outputs(4648));
    outputs(8762) <= layer2_outputs(10098);
    outputs(8763) <= (layer2_outputs(6850)) and (layer2_outputs(2746));
    outputs(8764) <= layer2_outputs(9930);
    outputs(8765) <= not(layer2_outputs(3553));
    outputs(8766) <= not(layer2_outputs(8296));
    outputs(8767) <= not(layer2_outputs(5749));
    outputs(8768) <= not((layer2_outputs(131)) or (layer2_outputs(9053)));
    outputs(8769) <= (layer2_outputs(5912)) and not (layer2_outputs(8474));
    outputs(8770) <= layer2_outputs(1706);
    outputs(8771) <= not(layer2_outputs(6413));
    outputs(8772) <= not((layer2_outputs(8573)) xor (layer2_outputs(7351)));
    outputs(8773) <= layer2_outputs(2146);
    outputs(8774) <= not(layer2_outputs(2689));
    outputs(8775) <= layer2_outputs(1871);
    outputs(8776) <= layer2_outputs(17);
    outputs(8777) <= layer2_outputs(1643);
    outputs(8778) <= (layer2_outputs(2402)) and not (layer2_outputs(5410));
    outputs(8779) <= layer2_outputs(9563);
    outputs(8780) <= layer2_outputs(5604);
    outputs(8781) <= layer2_outputs(4161);
    outputs(8782) <= not(layer2_outputs(3857));
    outputs(8783) <= not((layer2_outputs(3028)) or (layer2_outputs(3338)));
    outputs(8784) <= (layer2_outputs(7054)) xor (layer2_outputs(9185));
    outputs(8785) <= not(layer2_outputs(3581));
    outputs(8786) <= not(layer2_outputs(6296));
    outputs(8787) <= not(layer2_outputs(2492)) or (layer2_outputs(10135));
    outputs(8788) <= layer2_outputs(9032);
    outputs(8789) <= layer2_outputs(5686);
    outputs(8790) <= layer2_outputs(7045);
    outputs(8791) <= not((layer2_outputs(5364)) xor (layer2_outputs(8948)));
    outputs(8792) <= not(layer2_outputs(3845));
    outputs(8793) <= not((layer2_outputs(2287)) xor (layer2_outputs(5755)));
    outputs(8794) <= not(layer2_outputs(3904));
    outputs(8795) <= layer2_outputs(8028);
    outputs(8796) <= layer2_outputs(4229);
    outputs(8797) <= not((layer2_outputs(6100)) xor (layer2_outputs(3519)));
    outputs(8798) <= not(layer2_outputs(237));
    outputs(8799) <= not((layer2_outputs(6586)) xor (layer2_outputs(3832)));
    outputs(8800) <= not(layer2_outputs(7690));
    outputs(8801) <= layer2_outputs(5470);
    outputs(8802) <= not(layer2_outputs(1585));
    outputs(8803) <= not(layer2_outputs(9544));
    outputs(8804) <= not(layer2_outputs(1526));
    outputs(8805) <= not(layer2_outputs(7374));
    outputs(8806) <= layer2_outputs(2220);
    outputs(8807) <= not(layer2_outputs(361)) or (layer2_outputs(7673));
    outputs(8808) <= not(layer2_outputs(1561));
    outputs(8809) <= not(layer2_outputs(3648));
    outputs(8810) <= layer2_outputs(1352);
    outputs(8811) <= not(layer2_outputs(5978));
    outputs(8812) <= (layer2_outputs(8284)) or (layer2_outputs(9236));
    outputs(8813) <= (layer2_outputs(5442)) xor (layer2_outputs(2797));
    outputs(8814) <= not(layer2_outputs(8496));
    outputs(8815) <= layer2_outputs(4452);
    outputs(8816) <= not(layer2_outputs(1644));
    outputs(8817) <= (layer2_outputs(1653)) and (layer2_outputs(3693));
    outputs(8818) <= not((layer2_outputs(1630)) xor (layer2_outputs(6769)));
    outputs(8819) <= layer2_outputs(8710);
    outputs(8820) <= not((layer2_outputs(5847)) and (layer2_outputs(6037)));
    outputs(8821) <= (layer2_outputs(9640)) xor (layer2_outputs(4439));
    outputs(8822) <= not(layer2_outputs(2078));
    outputs(8823) <= not(layer2_outputs(9233));
    outputs(8824) <= not(layer2_outputs(6957));
    outputs(8825) <= not((layer2_outputs(8522)) xor (layer2_outputs(4970)));
    outputs(8826) <= not((layer2_outputs(6839)) xor (layer2_outputs(9419)));
    outputs(8827) <= layer2_outputs(4303);
    outputs(8828) <= not(layer2_outputs(4698));
    outputs(8829) <= (layer2_outputs(8559)) and not (layer2_outputs(2926));
    outputs(8830) <= not((layer2_outputs(5879)) xor (layer2_outputs(3424)));
    outputs(8831) <= not(layer2_outputs(4379)) or (layer2_outputs(1559));
    outputs(8832) <= not((layer2_outputs(8611)) and (layer2_outputs(9252)));
    outputs(8833) <= not((layer2_outputs(9269)) xor (layer2_outputs(2496)));
    outputs(8834) <= not(layer2_outputs(5229)) or (layer2_outputs(8400));
    outputs(8835) <= layer2_outputs(7681);
    outputs(8836) <= not(layer2_outputs(10057));
    outputs(8837) <= layer2_outputs(7181);
    outputs(8838) <= (layer2_outputs(5417)) and not (layer2_outputs(6304));
    outputs(8839) <= not(layer2_outputs(898)) or (layer2_outputs(973));
    outputs(8840) <= not(layer2_outputs(1283));
    outputs(8841) <= not((layer2_outputs(9496)) xor (layer2_outputs(687)));
    outputs(8842) <= not(layer2_outputs(1988));
    outputs(8843) <= layer2_outputs(9684);
    outputs(8844) <= not(layer2_outputs(8690));
    outputs(8845) <= (layer2_outputs(5387)) xor (layer2_outputs(6527));
    outputs(8846) <= (layer2_outputs(7733)) and not (layer2_outputs(6657));
    outputs(8847) <= (layer2_outputs(4862)) or (layer2_outputs(448));
    outputs(8848) <= (layer2_outputs(3267)) or (layer2_outputs(6052));
    outputs(8849) <= not(layer2_outputs(1367));
    outputs(8850) <= not((layer2_outputs(9874)) xor (layer2_outputs(9550)));
    outputs(8851) <= not((layer2_outputs(3703)) xor (layer2_outputs(7501)));
    outputs(8852) <= (layer2_outputs(4948)) xor (layer2_outputs(4334));
    outputs(8853) <= (layer2_outputs(2493)) xor (layer2_outputs(8263));
    outputs(8854) <= not(layer2_outputs(8007));
    outputs(8855) <= not(layer2_outputs(8557));
    outputs(8856) <= layer2_outputs(238);
    outputs(8857) <= not((layer2_outputs(5443)) xor (layer2_outputs(4430)));
    outputs(8858) <= (layer2_outputs(1588)) xor (layer2_outputs(8267));
    outputs(8859) <= layer2_outputs(519);
    outputs(8860) <= not((layer2_outputs(8980)) and (layer2_outputs(5635)));
    outputs(8861) <= not(layer2_outputs(10082)) or (layer2_outputs(9667));
    outputs(8862) <= not(layer2_outputs(6973));
    outputs(8863) <= (layer2_outputs(5778)) or (layer2_outputs(9826));
    outputs(8864) <= not((layer2_outputs(4868)) xor (layer2_outputs(2028)));
    outputs(8865) <= (layer2_outputs(8305)) xor (layer2_outputs(5077));
    outputs(8866) <= not((layer2_outputs(3412)) xor (layer2_outputs(8356)));
    outputs(8867) <= not((layer2_outputs(3417)) and (layer2_outputs(9141)));
    outputs(8868) <= (layer2_outputs(3138)) xor (layer2_outputs(7565));
    outputs(8869) <= (layer2_outputs(7830)) and not (layer2_outputs(4060));
    outputs(8870) <= layer2_outputs(6597);
    outputs(8871) <= not((layer2_outputs(4625)) or (layer2_outputs(4378)));
    outputs(8872) <= not((layer2_outputs(10174)) and (layer2_outputs(2753)));
    outputs(8873) <= (layer2_outputs(9855)) or (layer2_outputs(5880));
    outputs(8874) <= layer2_outputs(494);
    outputs(8875) <= not(layer2_outputs(8094)) or (layer2_outputs(7463));
    outputs(8876) <= not((layer2_outputs(9945)) xor (layer2_outputs(6726)));
    outputs(8877) <= not((layer2_outputs(3002)) and (layer2_outputs(247)));
    outputs(8878) <= not((layer2_outputs(4415)) xor (layer2_outputs(8278)));
    outputs(8879) <= (layer2_outputs(9852)) xor (layer2_outputs(6793));
    outputs(8880) <= not(layer2_outputs(1311));
    outputs(8881) <= (layer2_outputs(5042)) and not (layer2_outputs(7597));
    outputs(8882) <= layer2_outputs(3010);
    outputs(8883) <= (layer2_outputs(4320)) and not (layer2_outputs(1732));
    outputs(8884) <= not(layer2_outputs(4491)) or (layer2_outputs(7370));
    outputs(8885) <= not(layer2_outputs(7757));
    outputs(8886) <= layer2_outputs(5137);
    outputs(8887) <= not(layer2_outputs(858));
    outputs(8888) <= (layer2_outputs(9860)) xor (layer2_outputs(7745));
    outputs(8889) <= layer2_outputs(294);
    outputs(8890) <= (layer2_outputs(9784)) xor (layer2_outputs(2003));
    outputs(8891) <= not(layer2_outputs(7968)) or (layer2_outputs(8340));
    outputs(8892) <= not((layer2_outputs(8443)) and (layer2_outputs(1173)));
    outputs(8893) <= not((layer2_outputs(3453)) xor (layer2_outputs(4031)));
    outputs(8894) <= layer2_outputs(5980);
    outputs(8895) <= layer2_outputs(7700);
    outputs(8896) <= layer2_outputs(9460);
    outputs(8897) <= not((layer2_outputs(297)) xor (layer2_outputs(7049)));
    outputs(8898) <= not((layer2_outputs(5271)) and (layer2_outputs(4807)));
    outputs(8899) <= layer2_outputs(6770);
    outputs(8900) <= layer2_outputs(8393);
    outputs(8901) <= not(layer2_outputs(8725));
    outputs(8902) <= (layer2_outputs(895)) xor (layer2_outputs(3775));
    outputs(8903) <= not(layer2_outputs(3558));
    outputs(8904) <= not((layer2_outputs(4667)) xor (layer2_outputs(7359)));
    outputs(8905) <= layer2_outputs(3824);
    outputs(8906) <= not(layer2_outputs(4265));
    outputs(8907) <= not((layer2_outputs(10036)) xor (layer2_outputs(6334)));
    outputs(8908) <= layer2_outputs(8055);
    outputs(8909) <= (layer2_outputs(305)) and not (layer2_outputs(6470));
    outputs(8910) <= not((layer2_outputs(7833)) xor (layer2_outputs(5743)));
    outputs(8911) <= (layer2_outputs(4330)) xor (layer2_outputs(1032));
    outputs(8912) <= not((layer2_outputs(6071)) xor (layer2_outputs(9868)));
    outputs(8913) <= not(layer2_outputs(3661));
    outputs(8914) <= not((layer2_outputs(1567)) xor (layer2_outputs(8315)));
    outputs(8915) <= layer2_outputs(3974);
    outputs(8916) <= layer2_outputs(5794);
    outputs(8917) <= (layer2_outputs(1202)) xor (layer2_outputs(6187));
    outputs(8918) <= (layer2_outputs(6207)) xor (layer2_outputs(4558));
    outputs(8919) <= (layer2_outputs(3819)) and (layer2_outputs(505));
    outputs(8920) <= not((layer2_outputs(2726)) or (layer2_outputs(2364)));
    outputs(8921) <= not((layer2_outputs(7800)) xor (layer2_outputs(9359)));
    outputs(8922) <= not((layer2_outputs(7276)) xor (layer2_outputs(568)));
    outputs(8923) <= not((layer2_outputs(6094)) xor (layer2_outputs(1556)));
    outputs(8924) <= not(layer2_outputs(8730));
    outputs(8925) <= layer2_outputs(7775);
    outputs(8926) <= not(layer2_outputs(8703)) or (layer2_outputs(272));
    outputs(8927) <= (layer2_outputs(5105)) xor (layer2_outputs(5350));
    outputs(8928) <= not(layer2_outputs(2849));
    outputs(8929) <= not((layer2_outputs(9043)) xor (layer2_outputs(7514)));
    outputs(8930) <= not(layer2_outputs(452));
    outputs(8931) <= layer2_outputs(3466);
    outputs(8932) <= layer2_outputs(6027);
    outputs(8933) <= not((layer2_outputs(9984)) and (layer2_outputs(4276)));
    outputs(8934) <= not((layer2_outputs(6174)) xor (layer2_outputs(6694)));
    outputs(8935) <= not(layer2_outputs(1813));
    outputs(8936) <= not((layer2_outputs(10024)) xor (layer2_outputs(738)));
    outputs(8937) <= not(layer2_outputs(7252)) or (layer2_outputs(5396));
    outputs(8938) <= not(layer2_outputs(720));
    outputs(8939) <= not(layer2_outputs(4201));
    outputs(8940) <= layer2_outputs(6914);
    outputs(8941) <= not((layer2_outputs(757)) xor (layer2_outputs(7547)));
    outputs(8942) <= not(layer2_outputs(2213)) or (layer2_outputs(6585));
    outputs(8943) <= not(layer2_outputs(3762));
    outputs(8944) <= not((layer2_outputs(6457)) and (layer2_outputs(540)));
    outputs(8945) <= not((layer2_outputs(7000)) xor (layer2_outputs(9629)));
    outputs(8946) <= not(layer2_outputs(1644));
    outputs(8947) <= (layer2_outputs(4467)) or (layer2_outputs(6664));
    outputs(8948) <= layer2_outputs(6170);
    outputs(8949) <= layer2_outputs(9118);
    outputs(8950) <= (layer2_outputs(9976)) xor (layer2_outputs(9079));
    outputs(8951) <= not(layer2_outputs(4022));
    outputs(8952) <= layer2_outputs(9762);
    outputs(8953) <= layer2_outputs(5466);
    outputs(8954) <= not(layer2_outputs(3248));
    outputs(8955) <= not(layer2_outputs(9429)) or (layer2_outputs(9706));
    outputs(8956) <= not(layer2_outputs(2039));
    outputs(8957) <= not((layer2_outputs(1636)) and (layer2_outputs(3656)));
    outputs(8958) <= not(layer2_outputs(6509));
    outputs(8959) <= (layer2_outputs(4932)) xor (layer2_outputs(1836));
    outputs(8960) <= (layer2_outputs(6994)) and not (layer2_outputs(205));
    outputs(8961) <= not(layer2_outputs(8398));
    outputs(8962) <= not((layer2_outputs(5311)) xor (layer2_outputs(7577)));
    outputs(8963) <= (layer2_outputs(8874)) or (layer2_outputs(8820));
    outputs(8964) <= not((layer2_outputs(9037)) xor (layer2_outputs(132)));
    outputs(8965) <= not((layer2_outputs(6300)) and (layer2_outputs(9172)));
    outputs(8966) <= not(layer2_outputs(6350));
    outputs(8967) <= layer2_outputs(4693);
    outputs(8968) <= not((layer2_outputs(4059)) xor (layer2_outputs(9347)));
    outputs(8969) <= not((layer2_outputs(8105)) or (layer2_outputs(8372)));
    outputs(8970) <= layer2_outputs(7191);
    outputs(8971) <= not(layer2_outputs(5541));
    outputs(8972) <= not((layer2_outputs(9928)) xor (layer2_outputs(8719)));
    outputs(8973) <= layer2_outputs(4356);
    outputs(8974) <= (layer2_outputs(5530)) and not (layer2_outputs(1354));
    outputs(8975) <= (layer2_outputs(571)) xor (layer2_outputs(3136));
    outputs(8976) <= not(layer2_outputs(851));
    outputs(8977) <= not(layer2_outputs(4363)) or (layer2_outputs(8871));
    outputs(8978) <= (layer2_outputs(6416)) or (layer2_outputs(6478));
    outputs(8979) <= layer2_outputs(6830);
    outputs(8980) <= not(layer2_outputs(5662));
    outputs(8981) <= (layer2_outputs(10092)) xor (layer2_outputs(5909));
    outputs(8982) <= not(layer2_outputs(1638));
    outputs(8983) <= not(layer2_outputs(6526));
    outputs(8984) <= (layer2_outputs(2638)) xor (layer2_outputs(5679));
    outputs(8985) <= (layer2_outputs(2845)) or (layer2_outputs(4175));
    outputs(8986) <= not(layer2_outputs(1437)) or (layer2_outputs(801));
    outputs(8987) <= layer2_outputs(9276);
    outputs(8988) <= (layer2_outputs(5063)) xor (layer2_outputs(4027));
    outputs(8989) <= (layer2_outputs(5925)) xor (layer2_outputs(5391));
    outputs(8990) <= layer2_outputs(8547);
    outputs(8991) <= not((layer2_outputs(8420)) xor (layer2_outputs(146)));
    outputs(8992) <= not(layer2_outputs(3334)) or (layer2_outputs(3854));
    outputs(8993) <= (layer2_outputs(7855)) xor (layer2_outputs(4366));
    outputs(8994) <= not(layer2_outputs(8845));
    outputs(8995) <= not(layer2_outputs(3105));
    outputs(8996) <= layer2_outputs(1570);
    outputs(8997) <= not((layer2_outputs(4069)) xor (layer2_outputs(2141)));
    outputs(8998) <= (layer2_outputs(592)) xor (layer2_outputs(6796));
    outputs(8999) <= not(layer2_outputs(956));
    outputs(9000) <= not(layer2_outputs(224));
    outputs(9001) <= not((layer2_outputs(8011)) xor (layer2_outputs(6512)));
    outputs(9002) <= (layer2_outputs(7346)) xor (layer2_outputs(9435));
    outputs(9003) <= not(layer2_outputs(8624));
    outputs(9004) <= (layer2_outputs(6562)) xor (layer2_outputs(2023));
    outputs(9005) <= layer2_outputs(9607);
    outputs(9006) <= not((layer2_outputs(9130)) xor (layer2_outputs(7962)));
    outputs(9007) <= not(layer2_outputs(5863));
    outputs(9008) <= (layer2_outputs(2930)) or (layer2_outputs(4946));
    outputs(9009) <= not(layer2_outputs(9735));
    outputs(9010) <= not((layer2_outputs(1341)) xor (layer2_outputs(5578)));
    outputs(9011) <= not(layer2_outputs(1764)) or (layer2_outputs(4652));
    outputs(9012) <= not(layer2_outputs(9712));
    outputs(9013) <= not((layer2_outputs(6803)) xor (layer2_outputs(3010)));
    outputs(9014) <= layer2_outputs(2568);
    outputs(9015) <= not((layer2_outputs(1266)) xor (layer2_outputs(5035)));
    outputs(9016) <= not(layer2_outputs(3876));
    outputs(9017) <= not((layer2_outputs(10045)) xor (layer2_outputs(5438)));
    outputs(9018) <= not((layer2_outputs(308)) and (layer2_outputs(9737)));
    outputs(9019) <= not(layer2_outputs(963)) or (layer2_outputs(4293));
    outputs(9020) <= layer2_outputs(7914);
    outputs(9021) <= not((layer2_outputs(522)) xor (layer2_outputs(8109)));
    outputs(9022) <= (layer2_outputs(6277)) xor (layer2_outputs(6954));
    outputs(9023) <= (layer2_outputs(8021)) xor (layer2_outputs(9734));
    outputs(9024) <= (layer2_outputs(4964)) and (layer2_outputs(4888));
    outputs(9025) <= not(layer2_outputs(8069));
    outputs(9026) <= (layer2_outputs(5867)) or (layer2_outputs(396));
    outputs(9027) <= (layer2_outputs(3340)) and not (layer2_outputs(1627));
    outputs(9028) <= (layer2_outputs(6724)) xor (layer2_outputs(8765));
    outputs(9029) <= not(layer2_outputs(6532));
    outputs(9030) <= not(layer2_outputs(5516));
    outputs(9031) <= (layer2_outputs(5923)) xor (layer2_outputs(4515));
    outputs(9032) <= layer2_outputs(7347);
    outputs(9033) <= layer2_outputs(3478);
    outputs(9034) <= not(layer2_outputs(6647));
    outputs(9035) <= not(layer2_outputs(8096));
    outputs(9036) <= not((layer2_outputs(3978)) xor (layer2_outputs(6642)));
    outputs(9037) <= not((layer2_outputs(3842)) xor (layer2_outputs(6389)));
    outputs(9038) <= not(layer2_outputs(5623)) or (layer2_outputs(7202));
    outputs(9039) <= not(layer2_outputs(3352));
    outputs(9040) <= not((layer2_outputs(5312)) xor (layer2_outputs(9938)));
    outputs(9041) <= layer2_outputs(9824);
    outputs(9042) <= not((layer2_outputs(7376)) and (layer2_outputs(8909)));
    outputs(9043) <= not(layer2_outputs(4866)) or (layer2_outputs(8221));
    outputs(9044) <= (layer2_outputs(7685)) xor (layer2_outputs(9363));
    outputs(9045) <= (layer2_outputs(5002)) xor (layer2_outputs(7196));
    outputs(9046) <= not(layer2_outputs(5701));
    outputs(9047) <= layer2_outputs(3250);
    outputs(9048) <= not(layer2_outputs(3162));
    outputs(9049) <= (layer2_outputs(9364)) or (layer2_outputs(5112));
    outputs(9050) <= not(layer2_outputs(5617));
    outputs(9051) <= (layer2_outputs(2097)) xor (layer2_outputs(4527));
    outputs(9052) <= (layer2_outputs(3116)) xor (layer2_outputs(6166));
    outputs(9053) <= not(layer2_outputs(7317));
    outputs(9054) <= layer2_outputs(4623);
    outputs(9055) <= not(layer2_outputs(5126));
    outputs(9056) <= not((layer2_outputs(978)) xor (layer2_outputs(9859)));
    outputs(9057) <= not((layer2_outputs(6701)) xor (layer2_outputs(9201)));
    outputs(9058) <= not((layer2_outputs(5416)) xor (layer2_outputs(3275)));
    outputs(9059) <= layer2_outputs(9588);
    outputs(9060) <= layer2_outputs(9232);
    outputs(9061) <= not((layer2_outputs(4207)) xor (layer2_outputs(5531)));
    outputs(9062) <= (layer2_outputs(5165)) xor (layer2_outputs(4771));
    outputs(9063) <= (layer2_outputs(8382)) xor (layer2_outputs(3121));
    outputs(9064) <= (layer2_outputs(1322)) xor (layer2_outputs(3467));
    outputs(9065) <= not((layer2_outputs(855)) xor (layer2_outputs(1617)));
    outputs(9066) <= not((layer2_outputs(10099)) xor (layer2_outputs(9697)));
    outputs(9067) <= not(layer2_outputs(5556));
    outputs(9068) <= not((layer2_outputs(2628)) xor (layer2_outputs(6139)));
    outputs(9069) <= not((layer2_outputs(6199)) or (layer2_outputs(4779)));
    outputs(9070) <= layer2_outputs(3848);
    outputs(9071) <= not(layer2_outputs(4124));
    outputs(9072) <= not(layer2_outputs(9908)) or (layer2_outputs(8130));
    outputs(9073) <= not((layer2_outputs(4023)) and (layer2_outputs(2776)));
    outputs(9074) <= (layer2_outputs(3579)) xor (layer2_outputs(558));
    outputs(9075) <= not((layer2_outputs(9881)) xor (layer2_outputs(9160)));
    outputs(9076) <= not(layer2_outputs(4908));
    outputs(9077) <= layer2_outputs(487);
    outputs(9078) <= not(layer2_outputs(4400));
    outputs(9079) <= not(layer2_outputs(9046));
    outputs(9080) <= (layer2_outputs(2920)) xor (layer2_outputs(9711));
    outputs(9081) <= layer2_outputs(606);
    outputs(9082) <= (layer2_outputs(7824)) xor (layer2_outputs(139));
    outputs(9083) <= not((layer2_outputs(5995)) xor (layer2_outputs(6851)));
    outputs(9084) <= not((layer2_outputs(4296)) xor (layer2_outputs(1173)));
    outputs(9085) <= layer2_outputs(444);
    outputs(9086) <= layer2_outputs(5915);
    outputs(9087) <= not(layer2_outputs(7818));
    outputs(9088) <= not(layer2_outputs(25));
    outputs(9089) <= layer2_outputs(3274);
    outputs(9090) <= layer2_outputs(9214);
    outputs(9091) <= layer2_outputs(6063);
    outputs(9092) <= (layer2_outputs(9831)) and not (layer2_outputs(7818));
    outputs(9093) <= (layer2_outputs(4417)) xor (layer2_outputs(4173));
    outputs(9094) <= (layer2_outputs(6746)) and not (layer2_outputs(8205));
    outputs(9095) <= not((layer2_outputs(8566)) xor (layer2_outputs(1530)));
    outputs(9096) <= not(layer2_outputs(1184));
    outputs(9097) <= not(layer2_outputs(2684));
    outputs(9098) <= not((layer2_outputs(4040)) xor (layer2_outputs(8201)));
    outputs(9099) <= not(layer2_outputs(3415)) or (layer2_outputs(9527));
    outputs(9100) <= not((layer2_outputs(7028)) xor (layer2_outputs(2536)));
    outputs(9101) <= not((layer2_outputs(8405)) and (layer2_outputs(5973)));
    outputs(9102) <= not((layer2_outputs(8399)) xor (layer2_outputs(4070)));
    outputs(9103) <= (layer2_outputs(6051)) xor (layer2_outputs(4553));
    outputs(9104) <= not((layer2_outputs(9511)) xor (layer2_outputs(5513)));
    outputs(9105) <= not((layer2_outputs(317)) and (layer2_outputs(1497)));
    outputs(9106) <= (layer2_outputs(3113)) xor (layer2_outputs(3180));
    outputs(9107) <= layer2_outputs(7187);
    outputs(9108) <= layer2_outputs(1053);
    outputs(9109) <= layer2_outputs(8692);
    outputs(9110) <= not((layer2_outputs(8020)) xor (layer2_outputs(819)));
    outputs(9111) <= not((layer2_outputs(1821)) xor (layer2_outputs(2467)));
    outputs(9112) <= layer2_outputs(6682);
    outputs(9113) <= layer2_outputs(3481);
    outputs(9114) <= not((layer2_outputs(8705)) xor (layer2_outputs(1676)));
    outputs(9115) <= (layer2_outputs(7802)) xor (layer2_outputs(8810));
    outputs(9116) <= not((layer2_outputs(9851)) xor (layer2_outputs(8390)));
    outputs(9117) <= layer2_outputs(3708);
    outputs(9118) <= layer2_outputs(3922);
    outputs(9119) <= not(layer2_outputs(6934));
    outputs(9120) <= (layer2_outputs(8162)) or (layer2_outputs(5422));
    outputs(9121) <= layer2_outputs(658);
    outputs(9122) <= layer2_outputs(2063);
    outputs(9123) <= layer2_outputs(7274);
    outputs(9124) <= layer2_outputs(6287);
    outputs(9125) <= not(layer2_outputs(8008));
    outputs(9126) <= layer2_outputs(10181);
    outputs(9127) <= (layer2_outputs(9036)) xor (layer2_outputs(2310));
    outputs(9128) <= (layer2_outputs(265)) xor (layer2_outputs(5678));
    outputs(9129) <= not((layer2_outputs(1071)) and (layer2_outputs(2471)));
    outputs(9130) <= not((layer2_outputs(7285)) xor (layer2_outputs(2805)));
    outputs(9131) <= layer2_outputs(607);
    outputs(9132) <= not((layer2_outputs(6377)) xor (layer2_outputs(10103)));
    outputs(9133) <= not(layer2_outputs(6140));
    outputs(9134) <= layer2_outputs(4602);
    outputs(9135) <= layer2_outputs(1444);
    outputs(9136) <= not(layer2_outputs(7143));
    outputs(9137) <= layer2_outputs(8864);
    outputs(9138) <= not(layer2_outputs(2690));
    outputs(9139) <= not(layer2_outputs(1605)) or (layer2_outputs(7353));
    outputs(9140) <= (layer2_outputs(8815)) xor (layer2_outputs(2806));
    outputs(9141) <= not(layer2_outputs(7308)) or (layer2_outputs(3160));
    outputs(9142) <= not(layer2_outputs(6998));
    outputs(9143) <= not(layer2_outputs(821));
    outputs(9144) <= not(layer2_outputs(5620));
    outputs(9145) <= (layer2_outputs(3613)) xor (layer2_outputs(7751));
    outputs(9146) <= layer2_outputs(4075);
    outputs(9147) <= layer2_outputs(4639);
    outputs(9148) <= layer2_outputs(9309);
    outputs(9149) <= not(layer2_outputs(3403));
    outputs(9150) <= layer2_outputs(9167);
    outputs(9151) <= not((layer2_outputs(9396)) xor (layer2_outputs(4865)));
    outputs(9152) <= layer2_outputs(10204);
    outputs(9153) <= not(layer2_outputs(8139));
    outputs(9154) <= not((layer2_outputs(6780)) xor (layer2_outputs(8349)));
    outputs(9155) <= layer2_outputs(8898);
    outputs(9156) <= not((layer2_outputs(266)) xor (layer2_outputs(6800)));
    outputs(9157) <= layer2_outputs(2000);
    outputs(9158) <= not(layer2_outputs(4389));
    outputs(9159) <= not(layer2_outputs(3414));
    outputs(9160) <= not((layer2_outputs(6764)) xor (layer2_outputs(2544)));
    outputs(9161) <= layer2_outputs(3015);
    outputs(9162) <= layer2_outputs(5667);
    outputs(9163) <= not((layer2_outputs(5977)) and (layer2_outputs(3043)));
    outputs(9164) <= layer2_outputs(8402);
    outputs(9165) <= not((layer2_outputs(107)) xor (layer2_outputs(9145)));
    outputs(9166) <= layer2_outputs(7960);
    outputs(9167) <= layer2_outputs(1264);
    outputs(9168) <= not((layer2_outputs(2590)) xor (layer2_outputs(8968)));
    outputs(9169) <= (layer2_outputs(5299)) or (layer2_outputs(8841));
    outputs(9170) <= layer2_outputs(4135);
    outputs(9171) <= layer2_outputs(827);
    outputs(9172) <= layer2_outputs(6178);
    outputs(9173) <= not(layer2_outputs(4619));
    outputs(9174) <= not(layer2_outputs(7556));
    outputs(9175) <= (layer2_outputs(7767)) and not (layer2_outputs(9583));
    outputs(9176) <= layer2_outputs(10194);
    outputs(9177) <= (layer2_outputs(4335)) or (layer2_outputs(3951));
    outputs(9178) <= layer2_outputs(612);
    outputs(9179) <= not((layer2_outputs(5356)) xor (layer2_outputs(3391)));
    outputs(9180) <= layer2_outputs(3890);
    outputs(9181) <= layer2_outputs(6682);
    outputs(9182) <= layer2_outputs(3474);
    outputs(9183) <= not(layer2_outputs(7300));
    outputs(9184) <= not(layer2_outputs(8616));
    outputs(9185) <= not(layer2_outputs(9186));
    outputs(9186) <= (layer2_outputs(4391)) xor (layer2_outputs(6155));
    outputs(9187) <= layer2_outputs(8618);
    outputs(9188) <= not((layer2_outputs(4968)) xor (layer2_outputs(7212)));
    outputs(9189) <= not((layer2_outputs(3570)) xor (layer2_outputs(4854)));
    outputs(9190) <= not((layer2_outputs(5141)) xor (layer2_outputs(7643)));
    outputs(9191) <= not(layer2_outputs(919));
    outputs(9192) <= (layer2_outputs(180)) xor (layer2_outputs(339));
    outputs(9193) <= not(layer2_outputs(3987));
    outputs(9194) <= not((layer2_outputs(1422)) xor (layer2_outputs(9148)));
    outputs(9195) <= not((layer2_outputs(718)) xor (layer2_outputs(6898)));
    outputs(9196) <= not(layer2_outputs(670));
    outputs(9197) <= not(layer2_outputs(4533));
    outputs(9198) <= (layer2_outputs(6362)) xor (layer2_outputs(2122));
    outputs(9199) <= (layer2_outputs(2200)) xor (layer2_outputs(7883));
    outputs(9200) <= not((layer2_outputs(6566)) xor (layer2_outputs(3692)));
    outputs(9201) <= (layer2_outputs(4052)) xor (layer2_outputs(4376));
    outputs(9202) <= (layer2_outputs(9180)) xor (layer2_outputs(10077));
    outputs(9203) <= not(layer2_outputs(5483));
    outputs(9204) <= not(layer2_outputs(1246));
    outputs(9205) <= layer2_outputs(1483);
    outputs(9206) <= layer2_outputs(3213);
    outputs(9207) <= (layer2_outputs(748)) xor (layer2_outputs(3363));
    outputs(9208) <= not(layer2_outputs(2752));
    outputs(9209) <= not(layer2_outputs(1307));
    outputs(9210) <= not(layer2_outputs(3523));
    outputs(9211) <= layer2_outputs(8732);
    outputs(9212) <= not((layer2_outputs(1120)) xor (layer2_outputs(9713)));
    outputs(9213) <= (layer2_outputs(5824)) xor (layer2_outputs(8504));
    outputs(9214) <= not((layer2_outputs(5236)) xor (layer2_outputs(1934)));
    outputs(9215) <= layer2_outputs(10071);
    outputs(9216) <= not((layer2_outputs(3736)) xor (layer2_outputs(1597)));
    outputs(9217) <= layer2_outputs(1346);
    outputs(9218) <= (layer2_outputs(437)) and not (layer2_outputs(1466));
    outputs(9219) <= not(layer2_outputs(7628));
    outputs(9220) <= (layer2_outputs(4780)) and not (layer2_outputs(4227));
    outputs(9221) <= (layer2_outputs(4297)) and not (layer2_outputs(689));
    outputs(9222) <= layer2_outputs(6048);
    outputs(9223) <= (layer2_outputs(3375)) and not (layer2_outputs(3766));
    outputs(9224) <= not(layer2_outputs(7467));
    outputs(9225) <= layer2_outputs(8152);
    outputs(9226) <= layer2_outputs(4351);
    outputs(9227) <= not(layer2_outputs(4578));
    outputs(9228) <= (layer2_outputs(1693)) and (layer2_outputs(2885));
    outputs(9229) <= not(layer2_outputs(387));
    outputs(9230) <= (layer2_outputs(8086)) and (layer2_outputs(5733));
    outputs(9231) <= layer2_outputs(7211);
    outputs(9232) <= (layer2_outputs(2197)) and not (layer2_outputs(1594));
    outputs(9233) <= (layer2_outputs(7563)) and (layer2_outputs(7254));
    outputs(9234) <= layer2_outputs(4032);
    outputs(9235) <= not(layer2_outputs(1144));
    outputs(9236) <= not(layer2_outputs(8534));
    outputs(9237) <= not((layer2_outputs(9379)) and (layer2_outputs(1660)));
    outputs(9238) <= (layer2_outputs(7)) and not (layer2_outputs(2502));
    outputs(9239) <= layer2_outputs(6319);
    outputs(9240) <= (layer2_outputs(5888)) and (layer2_outputs(7977));
    outputs(9241) <= (layer2_outputs(9625)) and not (layer2_outputs(9351));
    outputs(9242) <= layer2_outputs(1509);
    outputs(9243) <= not((layer2_outputs(5090)) xor (layer2_outputs(2475)));
    outputs(9244) <= not(layer2_outputs(7214));
    outputs(9245) <= not((layer2_outputs(1778)) or (layer2_outputs(6700)));
    outputs(9246) <= not(layer2_outputs(497));
    outputs(9247) <= layer2_outputs(8157);
    outputs(9248) <= layer2_outputs(168);
    outputs(9249) <= not((layer2_outputs(9501)) xor (layer2_outputs(936)));
    outputs(9250) <= not(layer2_outputs(690));
    outputs(9251) <= (layer2_outputs(6388)) xor (layer2_outputs(5364));
    outputs(9252) <= not((layer2_outputs(3101)) xor (layer2_outputs(3359)));
    outputs(9253) <= layer2_outputs(8803);
    outputs(9254) <= not(layer2_outputs(8065)) or (layer2_outputs(1065));
    outputs(9255) <= (layer2_outputs(3302)) xor (layer2_outputs(4477));
    outputs(9256) <= not(layer2_outputs(4692));
    outputs(9257) <= layer2_outputs(2518);
    outputs(9258) <= (layer2_outputs(5998)) and not (layer2_outputs(9905));
    outputs(9259) <= not(layer2_outputs(6514));
    outputs(9260) <= not(layer2_outputs(5889));
    outputs(9261) <= not((layer2_outputs(1511)) xor (layer2_outputs(9774)));
    outputs(9262) <= layer2_outputs(2381);
    outputs(9263) <= not(layer2_outputs(3911));
    outputs(9264) <= (layer2_outputs(3000)) and not (layer2_outputs(1218));
    outputs(9265) <= not((layer2_outputs(7128)) xor (layer2_outputs(5322)));
    outputs(9266) <= not(layer2_outputs(1663));
    outputs(9267) <= layer2_outputs(2356);
    outputs(9268) <= not(layer2_outputs(3421));
    outputs(9269) <= not(layer2_outputs(5393));
    outputs(9270) <= not(layer2_outputs(4200));
    outputs(9271) <= (layer2_outputs(3060)) xor (layer2_outputs(5800));
    outputs(9272) <= layer2_outputs(1151);
    outputs(9273) <= layer2_outputs(9317);
    outputs(9274) <= (layer2_outputs(227)) xor (layer2_outputs(7307));
    outputs(9275) <= (layer2_outputs(139)) and not (layer2_outputs(444));
    outputs(9276) <= layer2_outputs(9271);
    outputs(9277) <= layer2_outputs(6064);
    outputs(9278) <= (layer2_outputs(1859)) and not (layer2_outputs(236));
    outputs(9279) <= not(layer2_outputs(9670));
    outputs(9280) <= not((layer2_outputs(4551)) xor (layer2_outputs(2812)));
    outputs(9281) <= not(layer2_outputs(5775));
    outputs(9282) <= (layer2_outputs(8981)) xor (layer2_outputs(770));
    outputs(9283) <= (layer2_outputs(7447)) and not (layer2_outputs(3867));
    outputs(9284) <= (layer2_outputs(4613)) or (layer2_outputs(6632));
    outputs(9285) <= not(layer2_outputs(2534));
    outputs(9286) <= (layer2_outputs(8876)) or (layer2_outputs(2807));
    outputs(9287) <= not(layer2_outputs(5060));
    outputs(9288) <= not(layer2_outputs(6568));
    outputs(9289) <= not((layer2_outputs(7788)) xor (layer2_outputs(4278)));
    outputs(9290) <= not(layer2_outputs(1520));
    outputs(9291) <= not(layer2_outputs(6098));
    outputs(9292) <= not((layer2_outputs(2997)) xor (layer2_outputs(6259)));
    outputs(9293) <= not(layer2_outputs(6741)) or (layer2_outputs(3065));
    outputs(9294) <= not(layer2_outputs(4458));
    outputs(9295) <= layer2_outputs(4435);
    outputs(9296) <= not((layer2_outputs(7159)) xor (layer2_outputs(6983)));
    outputs(9297) <= layer2_outputs(560);
    outputs(9298) <= layer2_outputs(6177);
    outputs(9299) <= not(layer2_outputs(4357));
    outputs(9300) <= not(layer2_outputs(8460));
    outputs(9301) <= (layer2_outputs(8278)) xor (layer2_outputs(10007));
    outputs(9302) <= layer2_outputs(1878);
    outputs(9303) <= (layer2_outputs(2446)) and (layer2_outputs(6751));
    outputs(9304) <= layer2_outputs(5862);
    outputs(9305) <= not((layer2_outputs(6744)) or (layer2_outputs(3656)));
    outputs(9306) <= layer2_outputs(835);
    outputs(9307) <= not(layer2_outputs(2182));
    outputs(9308) <= layer2_outputs(9533);
    outputs(9309) <= not(layer2_outputs(9925));
    outputs(9310) <= (layer2_outputs(1838)) and not (layer2_outputs(6624));
    outputs(9311) <= not(layer2_outputs(6882));
    outputs(9312) <= not(layer2_outputs(6876));
    outputs(9313) <= not(layer2_outputs(8916));
    outputs(9314) <= layer2_outputs(3365);
    outputs(9315) <= layer2_outputs(3108);
    outputs(9316) <= not(layer2_outputs(8995));
    outputs(9317) <= not(layer2_outputs(9033));
    outputs(9318) <= not(layer2_outputs(1253));
    outputs(9319) <= layer2_outputs(3050);
    outputs(9320) <= layer2_outputs(5004);
    outputs(9321) <= not(layer2_outputs(1098));
    outputs(9322) <= layer2_outputs(4716);
    outputs(9323) <= not((layer2_outputs(2439)) or (layer2_outputs(8004)));
    outputs(9324) <= (layer2_outputs(8760)) and (layer2_outputs(3527));
    outputs(9325) <= layer2_outputs(8297);
    outputs(9326) <= not(layer2_outputs(2231));
    outputs(9327) <= not((layer2_outputs(746)) or (layer2_outputs(7248)));
    outputs(9328) <= not(layer2_outputs(8984));
    outputs(9329) <= not(layer2_outputs(7545));
    outputs(9330) <= (layer2_outputs(8457)) xor (layer2_outputs(7995));
    outputs(9331) <= (layer2_outputs(2516)) or (layer2_outputs(4998));
    outputs(9332) <= not(layer2_outputs(7969)) or (layer2_outputs(9823));
    outputs(9333) <= layer2_outputs(5564);
    outputs(9334) <= (layer2_outputs(1633)) and not (layer2_outputs(3508));
    outputs(9335) <= (layer2_outputs(938)) or (layer2_outputs(4168));
    outputs(9336) <= layer2_outputs(7618);
    outputs(9337) <= (layer2_outputs(4383)) xor (layer2_outputs(2633));
    outputs(9338) <= not(layer2_outputs(8604));
    outputs(9339) <= not(layer2_outputs(2813));
    outputs(9340) <= layer2_outputs(613);
    outputs(9341) <= not(layer2_outputs(9050));
    outputs(9342) <= layer2_outputs(7297);
    outputs(9343) <= (layer2_outputs(2747)) and (layer2_outputs(8160));
    outputs(9344) <= not((layer2_outputs(7191)) xor (layer2_outputs(6015)));
    outputs(9345) <= layer2_outputs(6186);
    outputs(9346) <= not(layer2_outputs(2498)) or (layer2_outputs(3893));
    outputs(9347) <= not(layer2_outputs(6266)) or (layer2_outputs(8432));
    outputs(9348) <= layer2_outputs(6387);
    outputs(9349) <= (layer2_outputs(7928)) and not (layer2_outputs(1142));
    outputs(9350) <= (layer2_outputs(9962)) xor (layer2_outputs(1785));
    outputs(9351) <= not(layer2_outputs(5428));
    outputs(9352) <= layer2_outputs(9551);
    outputs(9353) <= not(layer2_outputs(772));
    outputs(9354) <= not((layer2_outputs(1564)) or (layer2_outputs(3096)));
    outputs(9355) <= (layer2_outputs(4961)) xor (layer2_outputs(7785));
    outputs(9356) <= not(layer2_outputs(1934));
    outputs(9357) <= layer2_outputs(1156);
    outputs(9358) <= not((layer2_outputs(1564)) xor (layer2_outputs(4089)));
    outputs(9359) <= (layer2_outputs(6649)) xor (layer2_outputs(8858));
    outputs(9360) <= not((layer2_outputs(5329)) xor (layer2_outputs(7533)));
    outputs(9361) <= layer2_outputs(6644);
    outputs(9362) <= not(layer2_outputs(397)) or (layer2_outputs(4094));
    outputs(9363) <= layer2_outputs(8159);
    outputs(9364) <= not((layer2_outputs(7674)) and (layer2_outputs(8079)));
    outputs(9365) <= layer2_outputs(7140);
    outputs(9366) <= not(layer2_outputs(1031));
    outputs(9367) <= not((layer2_outputs(4441)) xor (layer2_outputs(7571)));
    outputs(9368) <= (layer2_outputs(10085)) xor (layer2_outputs(7830));
    outputs(9369) <= not(layer2_outputs(2892));
    outputs(9370) <= not((layer2_outputs(4786)) or (layer2_outputs(9142)));
    outputs(9371) <= (layer2_outputs(7295)) xor (layer2_outputs(6084));
    outputs(9372) <= (layer2_outputs(6111)) and (layer2_outputs(8781));
    outputs(9373) <= not(layer2_outputs(7732));
    outputs(9374) <= (layer2_outputs(1140)) xor (layer2_outputs(10224));
    outputs(9375) <= layer2_outputs(137);
    outputs(9376) <= (layer2_outputs(5379)) xor (layer2_outputs(4488));
    outputs(9377) <= not(layer2_outputs(3266));
    outputs(9378) <= layer2_outputs(4586);
    outputs(9379) <= layer2_outputs(7314);
    outputs(9380) <= layer2_outputs(5702);
    outputs(9381) <= (layer2_outputs(9483)) and (layer2_outputs(288));
    outputs(9382) <= (layer2_outputs(2004)) and not (layer2_outputs(5270));
    outputs(9383) <= (layer2_outputs(6382)) and not (layer2_outputs(4026));
    outputs(9384) <= layer2_outputs(41);
    outputs(9385) <= not((layer2_outputs(3928)) xor (layer2_outputs(8238)));
    outputs(9386) <= not(layer2_outputs(8641)) or (layer2_outputs(2247));
    outputs(9387) <= (layer2_outputs(5513)) and not (layer2_outputs(8551));
    outputs(9388) <= not(layer2_outputs(3588));
    outputs(9389) <= layer2_outputs(7092);
    outputs(9390) <= not((layer2_outputs(2201)) xor (layer2_outputs(3088)));
    outputs(9391) <= not(layer2_outputs(3578));
    outputs(9392) <= not(layer2_outputs(4933));
    outputs(9393) <= (layer2_outputs(5401)) and not (layer2_outputs(7776));
    outputs(9394) <= not((layer2_outputs(3198)) xor (layer2_outputs(4551)));
    outputs(9395) <= not(layer2_outputs(1719));
    outputs(9396) <= not(layer2_outputs(7001));
    outputs(9397) <= (layer2_outputs(4264)) and not (layer2_outputs(405));
    outputs(9398) <= not(layer2_outputs(4483)) or (layer2_outputs(7923));
    outputs(9399) <= not(layer2_outputs(2134));
    outputs(9400) <= layer2_outputs(1943);
    outputs(9401) <= not(layer2_outputs(285));
    outputs(9402) <= (layer2_outputs(4677)) xor (layer2_outputs(5214));
    outputs(9403) <= not((layer2_outputs(8116)) and (layer2_outputs(3218)));
    outputs(9404) <= not(layer2_outputs(1506));
    outputs(9405) <= not((layer2_outputs(906)) or (layer2_outputs(5792)));
    outputs(9406) <= (layer2_outputs(2619)) and not (layer2_outputs(2231));
    outputs(9407) <= layer2_outputs(2661);
    outputs(9408) <= (layer2_outputs(4)) and (layer2_outputs(3411));
    outputs(9409) <= not((layer2_outputs(5103)) or (layer2_outputs(8879)));
    outputs(9410) <= (layer2_outputs(7687)) xor (layer2_outputs(4497));
    outputs(9411) <= (layer2_outputs(9235)) and (layer2_outputs(1767));
    outputs(9412) <= not(layer2_outputs(4538));
    outputs(9413) <= layer2_outputs(1174);
    outputs(9414) <= layer2_outputs(3162);
    outputs(9415) <= not((layer2_outputs(8372)) xor (layer2_outputs(1515)));
    outputs(9416) <= layer2_outputs(6716);
    outputs(9417) <= not(layer2_outputs(8895));
    outputs(9418) <= (layer2_outputs(6230)) and not (layer2_outputs(26));
    outputs(9419) <= (layer2_outputs(7023)) and (layer2_outputs(3716));
    outputs(9420) <= layer2_outputs(2306);
    outputs(9421) <= not((layer2_outputs(6422)) or (layer2_outputs(10084)));
    outputs(9422) <= not((layer2_outputs(4451)) xor (layer2_outputs(8247)));
    outputs(9423) <= not(layer2_outputs(6312));
    outputs(9424) <= not(layer2_outputs(3313));
    outputs(9425) <= not((layer2_outputs(5839)) xor (layer2_outputs(2798)));
    outputs(9426) <= layer2_outputs(7924);
    outputs(9427) <= (layer2_outputs(1807)) and not (layer2_outputs(6482));
    outputs(9428) <= (layer2_outputs(7238)) xor (layer2_outputs(1474));
    outputs(9429) <= (layer2_outputs(6520)) and not (layer2_outputs(1683));
    outputs(9430) <= not(layer2_outputs(8442));
    outputs(9431) <= (layer2_outputs(5506)) xor (layer2_outputs(5849));
    outputs(9432) <= not(layer2_outputs(1548));
    outputs(9433) <= not((layer2_outputs(3917)) xor (layer2_outputs(5526)));
    outputs(9434) <= (layer2_outputs(2032)) or (layer2_outputs(7234));
    outputs(9435) <= layer2_outputs(3531);
    outputs(9436) <= layer2_outputs(9528);
    outputs(9437) <= (layer2_outputs(9479)) and not (layer2_outputs(806));
    outputs(9438) <= not((layer2_outputs(8565)) xor (layer2_outputs(3688)));
    outputs(9439) <= not((layer2_outputs(5696)) or (layer2_outputs(218)));
    outputs(9440) <= (layer2_outputs(8695)) xor (layer2_outputs(10108));
    outputs(9441) <= layer2_outputs(5382);
    outputs(9442) <= layer2_outputs(1849);
    outputs(9443) <= not((layer2_outputs(839)) and (layer2_outputs(1635)));
    outputs(9444) <= (layer2_outputs(8525)) xor (layer2_outputs(4668));
    outputs(9445) <= not(layer2_outputs(7328));
    outputs(9446) <= not(layer2_outputs(5964));
    outputs(9447) <= not((layer2_outputs(2112)) xor (layer2_outputs(2737)));
    outputs(9448) <= layer2_outputs(4563);
    outputs(9449) <= not((layer2_outputs(3933)) or (layer2_outputs(7081)));
    outputs(9450) <= (layer2_outputs(1480)) and not (layer2_outputs(8117));
    outputs(9451) <= not(layer2_outputs(6693));
    outputs(9452) <= (layer2_outputs(4277)) xor (layer2_outputs(9972));
    outputs(9453) <= not(layer2_outputs(64));
    outputs(9454) <= not((layer2_outputs(4985)) and (layer2_outputs(4673)));
    outputs(9455) <= not(layer2_outputs(8720));
    outputs(9456) <= layer2_outputs(5266);
    outputs(9457) <= layer2_outputs(2405);
    outputs(9458) <= not(layer2_outputs(6997));
    outputs(9459) <= layer2_outputs(9292);
    outputs(9460) <= layer2_outputs(2374);
    outputs(9461) <= layer2_outputs(5063);
    outputs(9462) <= layer2_outputs(1546);
    outputs(9463) <= (layer2_outputs(2317)) xor (layer2_outputs(2850));
    outputs(9464) <= (layer2_outputs(1973)) and (layer2_outputs(9211));
    outputs(9465) <= not((layer2_outputs(9528)) xor (layer2_outputs(8668)));
    outputs(9466) <= (layer2_outputs(1205)) and not (layer2_outputs(7350));
    outputs(9467) <= layer2_outputs(9408);
    outputs(9468) <= layer2_outputs(9221);
    outputs(9469) <= (layer2_outputs(7881)) and not (layer2_outputs(1079));
    outputs(9470) <= layer2_outputs(590);
    outputs(9471) <= (layer2_outputs(8448)) xor (layer2_outputs(2145));
    outputs(9472) <= not(layer2_outputs(7287));
    outputs(9473) <= not(layer2_outputs(8388));
    outputs(9474) <= (layer2_outputs(101)) or (layer2_outputs(3889));
    outputs(9475) <= not(layer2_outputs(6318));
    outputs(9476) <= (layer2_outputs(295)) and not (layer2_outputs(2062));
    outputs(9477) <= not(layer2_outputs(7549));
    outputs(9478) <= not((layer2_outputs(3534)) xor (layer2_outputs(1070)));
    outputs(9479) <= (layer2_outputs(9102)) xor (layer2_outputs(2327));
    outputs(9480) <= layer2_outputs(6154);
    outputs(9481) <= not(layer2_outputs(7766));
    outputs(9482) <= (layer2_outputs(2322)) xor (layer2_outputs(5708));
    outputs(9483) <= not((layer2_outputs(7740)) xor (layer2_outputs(1842)));
    outputs(9484) <= layer2_outputs(3327);
    outputs(9485) <= layer2_outputs(8967);
    outputs(9486) <= not(layer2_outputs(4997));
    outputs(9487) <= (layer2_outputs(9062)) and not (layer2_outputs(3632));
    outputs(9488) <= not((layer2_outputs(9344)) xor (layer2_outputs(8261)));
    outputs(9489) <= layer2_outputs(3154);
    outputs(9490) <= layer2_outputs(2218);
    outputs(9491) <= not(layer2_outputs(3818));
    outputs(9492) <= not(layer2_outputs(7364));
    outputs(9493) <= (layer2_outputs(3387)) and not (layer2_outputs(2857));
    outputs(9494) <= not(layer2_outputs(1274));
    outputs(9495) <= not((layer2_outputs(1826)) and (layer2_outputs(6073)));
    outputs(9496) <= layer2_outputs(8482);
    outputs(9497) <= layer2_outputs(1895);
    outputs(9498) <= not(layer2_outputs(9547));
    outputs(9499) <= (layer2_outputs(1417)) and (layer2_outputs(4037));
    outputs(9500) <= not((layer2_outputs(1090)) xor (layer2_outputs(588)));
    outputs(9501) <= not(layer2_outputs(9814));
    outputs(9502) <= (layer2_outputs(8622)) and not (layer2_outputs(1286));
    outputs(9503) <= not(layer2_outputs(6805));
    outputs(9504) <= (layer2_outputs(2614)) and not (layer2_outputs(8290));
    outputs(9505) <= (layer2_outputs(7073)) and (layer2_outputs(5310));
    outputs(9506) <= layer2_outputs(376);
    outputs(9507) <= (layer2_outputs(6471)) or (layer2_outputs(6173));
    outputs(9508) <= layer2_outputs(4670);
    outputs(9509) <= layer2_outputs(5898);
    outputs(9510) <= not(layer2_outputs(1712));
    outputs(9511) <= (layer2_outputs(1904)) and not (layer2_outputs(1006));
    outputs(9512) <= layer2_outputs(4192);
    outputs(9513) <= not(layer2_outputs(584)) or (layer2_outputs(7102));
    outputs(9514) <= layer2_outputs(4157);
    outputs(9515) <= layer2_outputs(7620);
    outputs(9516) <= layer2_outputs(9342);
    outputs(9517) <= (layer2_outputs(5614)) or (layer2_outputs(5475));
    outputs(9518) <= (layer2_outputs(10097)) and (layer2_outputs(3710));
    outputs(9519) <= not((layer2_outputs(6910)) or (layer2_outputs(6191)));
    outputs(9520) <= layer2_outputs(2315);
    outputs(9521) <= (layer2_outputs(2387)) xor (layer2_outputs(9458));
    outputs(9522) <= layer2_outputs(5006);
    outputs(9523) <= layer2_outputs(1038);
    outputs(9524) <= not(layer2_outputs(2238));
    outputs(9525) <= layer2_outputs(2047);
    outputs(9526) <= not(layer2_outputs(9612));
    outputs(9527) <= not(layer2_outputs(3624));
    outputs(9528) <= (layer2_outputs(1886)) and not (layer2_outputs(2076));
    outputs(9529) <= not((layer2_outputs(6789)) or (layer2_outputs(6587)));
    outputs(9530) <= not((layer2_outputs(3605)) xor (layer2_outputs(4118)));
    outputs(9531) <= (layer2_outputs(5519)) xor (layer2_outputs(3790));
    outputs(9532) <= not((layer2_outputs(3770)) or (layer2_outputs(365)));
    outputs(9533) <= (layer2_outputs(378)) xor (layer2_outputs(8039));
    outputs(9534) <= not((layer2_outputs(6169)) xor (layer2_outputs(3774)));
    outputs(9535) <= (layer2_outputs(9212)) xor (layer2_outputs(2060));
    outputs(9536) <= not(layer2_outputs(2506));
    outputs(9537) <= not(layer2_outputs(711));
    outputs(9538) <= not(layer2_outputs(7979));
    outputs(9539) <= not((layer2_outputs(10160)) xor (layer2_outputs(6618)));
    outputs(9540) <= not(layer2_outputs(1783));
    outputs(9541) <= layer2_outputs(9451);
    outputs(9542) <= (layer2_outputs(8751)) and not (layer2_outputs(3471));
    outputs(9543) <= layer2_outputs(5385);
    outputs(9544) <= not(layer2_outputs(6005));
    outputs(9545) <= (layer2_outputs(6006)) xor (layer2_outputs(6945));
    outputs(9546) <= not(layer2_outputs(5158));
    outputs(9547) <= not(layer2_outputs(2418));
    outputs(9548) <= (layer2_outputs(4674)) xor (layer2_outputs(4912));
    outputs(9549) <= (layer2_outputs(7753)) xor (layer2_outputs(1863));
    outputs(9550) <= (layer2_outputs(5249)) and (layer2_outputs(9107));
    outputs(9551) <= layer2_outputs(9551);
    outputs(9552) <= layer2_outputs(2762);
    outputs(9553) <= not((layer2_outputs(2878)) xor (layer2_outputs(1395)));
    outputs(9554) <= layer2_outputs(1942);
    outputs(9555) <= layer2_outputs(1910);
    outputs(9556) <= not(layer2_outputs(5328));
    outputs(9557) <= not(layer2_outputs(3567));
    outputs(9558) <= not(layer2_outputs(1639));
    outputs(9559) <= not(layer2_outputs(4768));
    outputs(9560) <= not((layer2_outputs(10231)) xor (layer2_outputs(9466)));
    outputs(9561) <= layer2_outputs(2537);
    outputs(9562) <= not((layer2_outputs(8424)) xor (layer2_outputs(9783)));
    outputs(9563) <= not(layer2_outputs(2604));
    outputs(9564) <= not(layer2_outputs(6514));
    outputs(9565) <= not(layer2_outputs(9885));
    outputs(9566) <= not(layer2_outputs(1816));
    outputs(9567) <= not((layer2_outputs(6250)) xor (layer2_outputs(2355)));
    outputs(9568) <= not(layer2_outputs(702));
    outputs(9569) <= layer2_outputs(7332);
    outputs(9570) <= layer2_outputs(8554);
    outputs(9571) <= layer2_outputs(8463);
    outputs(9572) <= not(layer2_outputs(3617));
    outputs(9573) <= (layer2_outputs(5379)) and (layer2_outputs(399));
    outputs(9574) <= not((layer2_outputs(4749)) xor (layer2_outputs(6825)));
    outputs(9575) <= layer2_outputs(883);
    outputs(9576) <= layer2_outputs(7645);
    outputs(9577) <= layer2_outputs(4560);
    outputs(9578) <= not(layer2_outputs(6577)) or (layer2_outputs(6782));
    outputs(9579) <= layer2_outputs(8168);
    outputs(9580) <= (layer2_outputs(9537)) xor (layer2_outputs(3279));
    outputs(9581) <= layer2_outputs(6976);
    outputs(9582) <= (layer2_outputs(9639)) and (layer2_outputs(1713));
    outputs(9583) <= not(layer2_outputs(6574));
    outputs(9584) <= not(layer2_outputs(8585));
    outputs(9585) <= (layer2_outputs(3487)) and (layer2_outputs(8162));
    outputs(9586) <= not(layer2_outputs(4627));
    outputs(9587) <= (layer2_outputs(4672)) xor (layer2_outputs(779));
    outputs(9588) <= layer2_outputs(8358);
    outputs(9589) <= layer2_outputs(3853);
    outputs(9590) <= (layer2_outputs(10090)) and not (layer2_outputs(2900));
    outputs(9591) <= not(layer2_outputs(4566)) or (layer2_outputs(1531));
    outputs(9592) <= not(layer2_outputs(10077));
    outputs(9593) <= not(layer2_outputs(5316));
    outputs(9594) <= not(layer2_outputs(3374));
    outputs(9595) <= (layer2_outputs(9269)) or (layer2_outputs(9503));
    outputs(9596) <= not(layer2_outputs(9911));
    outputs(9597) <= (layer2_outputs(4870)) and (layer2_outputs(9147));
    outputs(9598) <= (layer2_outputs(9520)) and (layer2_outputs(9771));
    outputs(9599) <= not(layer2_outputs(6239));
    outputs(9600) <= not(layer2_outputs(760));
    outputs(9601) <= (layer2_outputs(6746)) xor (layer2_outputs(7136));
    outputs(9602) <= not(layer2_outputs(3169));
    outputs(9603) <= not((layer2_outputs(6951)) or (layer2_outputs(8195)));
    outputs(9604) <= not(layer2_outputs(4163));
    outputs(9605) <= not(layer2_outputs(5706));
    outputs(9606) <= (layer2_outputs(4036)) xor (layer2_outputs(1952));
    outputs(9607) <= not(layer2_outputs(4105));
    outputs(9608) <= (layer2_outputs(6018)) xor (layer2_outputs(5795));
    outputs(9609) <= layer2_outputs(168);
    outputs(9610) <= not(layer2_outputs(8370));
    outputs(9611) <= not(layer2_outputs(5872));
    outputs(9612) <= (layer2_outputs(4351)) and not (layer2_outputs(2756));
    outputs(9613) <= layer2_outputs(597);
    outputs(9614) <= not((layer2_outputs(6582)) and (layer2_outputs(1263)));
    outputs(9615) <= not(layer2_outputs(7506));
    outputs(9616) <= not(layer2_outputs(1952));
    outputs(9617) <= (layer2_outputs(1036)) or (layer2_outputs(3627));
    outputs(9618) <= not((layer2_outputs(5763)) and (layer2_outputs(6598)));
    outputs(9619) <= (layer2_outputs(3289)) or (layer2_outputs(7808));
    outputs(9620) <= not(layer2_outputs(1773));
    outputs(9621) <= not(layer2_outputs(8227));
    outputs(9622) <= (layer2_outputs(2475)) or (layer2_outputs(6112));
    outputs(9623) <= not(layer2_outputs(10062)) or (layer2_outputs(7420));
    outputs(9624) <= layer2_outputs(9462);
    outputs(9625) <= not(layer2_outputs(6448));
    outputs(9626) <= layer2_outputs(9196);
    outputs(9627) <= not(layer2_outputs(7994));
    outputs(9628) <= layer2_outputs(7083);
    outputs(9629) <= (layer2_outputs(7480)) or (layer2_outputs(341));
    outputs(9630) <= (layer2_outputs(6780)) xor (layer2_outputs(4869));
    outputs(9631) <= (layer2_outputs(1068)) and not (layer2_outputs(5881));
    outputs(9632) <= layer2_outputs(7941);
    outputs(9633) <= (layer2_outputs(8184)) or (layer2_outputs(6738));
    outputs(9634) <= not(layer2_outputs(6335));
    outputs(9635) <= layer2_outputs(1386);
    outputs(9636) <= not(layer2_outputs(2567)) or (layer2_outputs(4864));
    outputs(9637) <= not((layer2_outputs(4981)) or (layer2_outputs(9604)));
    outputs(9638) <= layer2_outputs(5424);
    outputs(9639) <= not(layer2_outputs(3252));
    outputs(9640) <= (layer2_outputs(3560)) xor (layer2_outputs(9621));
    outputs(9641) <= layer2_outputs(458);
    outputs(9642) <= not((layer2_outputs(7834)) xor (layer2_outputs(7779)));
    outputs(9643) <= not(layer2_outputs(6453));
    outputs(9644) <= layer2_outputs(1193);
    outputs(9645) <= (layer2_outputs(6678)) and not (layer2_outputs(2190));
    outputs(9646) <= (layer2_outputs(6706)) or (layer2_outputs(9778));
    outputs(9647) <= not(layer2_outputs(3639));
    outputs(9648) <= layer2_outputs(3027);
    outputs(9649) <= not(layer2_outputs(8704));
    outputs(9650) <= layer2_outputs(9728);
    outputs(9651) <= not(layer2_outputs(1683));
    outputs(9652) <= layer2_outputs(5068);
    outputs(9653) <= not(layer2_outputs(5720));
    outputs(9654) <= not(layer2_outputs(141));
    outputs(9655) <= (layer2_outputs(3956)) and not (layer2_outputs(5394));
    outputs(9656) <= not(layer2_outputs(8694));
    outputs(9657) <= (layer2_outputs(4574)) xor (layer2_outputs(76));
    outputs(9658) <= not(layer2_outputs(9356)) or (layer2_outputs(10004));
    outputs(9659) <= (layer2_outputs(3034)) xor (layer2_outputs(3446));
    outputs(9660) <= not((layer2_outputs(9864)) xor (layer2_outputs(39)));
    outputs(9661) <= (layer2_outputs(6676)) and (layer2_outputs(7631));
    outputs(9662) <= not((layer2_outputs(7406)) xor (layer2_outputs(1966)));
    outputs(9663) <= not(layer2_outputs(478));
    outputs(9664) <= not((layer2_outputs(10083)) xor (layer2_outputs(4946)));
    outputs(9665) <= layer2_outputs(766);
    outputs(9666) <= not(layer2_outputs(4587));
    outputs(9667) <= layer2_outputs(726);
    outputs(9668) <= (layer2_outputs(8164)) and not (layer2_outputs(9518));
    outputs(9669) <= (layer2_outputs(842)) xor (layer2_outputs(2887));
    outputs(9670) <= layer2_outputs(8794);
    outputs(9671) <= (layer2_outputs(95)) xor (layer2_outputs(1471));
    outputs(9672) <= not((layer2_outputs(3977)) xor (layer2_outputs(2565)));
    outputs(9673) <= layer2_outputs(3864);
    outputs(9674) <= (layer2_outputs(9948)) xor (layer2_outputs(7291));
    outputs(9675) <= layer2_outputs(10115);
    outputs(9676) <= (layer2_outputs(5098)) and (layer2_outputs(6921));
    outputs(9677) <= not(layer2_outputs(7156));
    outputs(9678) <= not(layer2_outputs(4481));
    outputs(9679) <= (layer2_outputs(8886)) and (layer2_outputs(2297));
    outputs(9680) <= layer2_outputs(3495);
    outputs(9681) <= not(layer2_outputs(4274));
    outputs(9682) <= (layer2_outputs(6496)) xor (layer2_outputs(6273));
    outputs(9683) <= layer2_outputs(2386);
    outputs(9684) <= (layer2_outputs(9647)) xor (layer2_outputs(273));
    outputs(9685) <= not(layer2_outputs(566)) or (layer2_outputs(4685));
    outputs(9686) <= (layer2_outputs(10088)) and not (layer2_outputs(4380));
    outputs(9687) <= (layer2_outputs(6504)) and not (layer2_outputs(7425));
    outputs(9688) <= (layer2_outputs(9395)) xor (layer2_outputs(3481));
    outputs(9689) <= (layer2_outputs(6446)) or (layer2_outputs(4052));
    outputs(9690) <= not(layer2_outputs(8784));
    outputs(9691) <= layer2_outputs(9643);
    outputs(9692) <= not(layer2_outputs(4852)) or (layer2_outputs(8331));
    outputs(9693) <= not(layer2_outputs(8585)) or (layer2_outputs(9386));
    outputs(9694) <= not(layer2_outputs(7015));
    outputs(9695) <= layer2_outputs(2870);
    outputs(9696) <= (layer2_outputs(7354)) and (layer2_outputs(9834));
    outputs(9697) <= not(layer2_outputs(7588));
    outputs(9698) <= layer2_outputs(230);
    outputs(9699) <= (layer2_outputs(6326)) xor (layer2_outputs(7039));
    outputs(9700) <= layer2_outputs(2645);
    outputs(9701) <= not(layer2_outputs(3583));
    outputs(9702) <= layer2_outputs(8363);
    outputs(9703) <= layer2_outputs(2601);
    outputs(9704) <= not(layer2_outputs(3268));
    outputs(9705) <= layer2_outputs(7434);
    outputs(9706) <= (layer2_outputs(6454)) and not (layer2_outputs(1557));
    outputs(9707) <= (layer2_outputs(6212)) and not (layer2_outputs(7060));
    outputs(9708) <= not((layer2_outputs(4195)) xor (layer2_outputs(115)));
    outputs(9709) <= layer2_outputs(5503);
    outputs(9710) <= not(layer2_outputs(7012));
    outputs(9711) <= not((layer2_outputs(4836)) xor (layer2_outputs(8687)));
    outputs(9712) <= not(layer2_outputs(7213));
    outputs(9713) <= (layer2_outputs(7082)) or (layer2_outputs(591));
    outputs(9714) <= not((layer2_outputs(2032)) xor (layer2_outputs(5500)));
    outputs(9715) <= not((layer2_outputs(2113)) or (layer2_outputs(9593)));
    outputs(9716) <= not(layer2_outputs(5107));
    outputs(9717) <= layer2_outputs(426);
    outputs(9718) <= not((layer2_outputs(181)) xor (layer2_outputs(110)));
    outputs(9719) <= not(layer2_outputs(5777));
    outputs(9720) <= (layer2_outputs(939)) and (layer2_outputs(5383));
    outputs(9721) <= (layer2_outputs(5949)) xor (layer2_outputs(6148));
    outputs(9722) <= (layer2_outputs(8158)) xor (layer2_outputs(6043));
    outputs(9723) <= not(layer2_outputs(5990));
    outputs(9724) <= not((layer2_outputs(8452)) and (layer2_outputs(1611)));
    outputs(9725) <= not(layer2_outputs(7034)) or (layer2_outputs(1078));
    outputs(9726) <= not(layer2_outputs(9));
    outputs(9727) <= (layer2_outputs(4207)) xor (layer2_outputs(8786));
    outputs(9728) <= layer2_outputs(2246);
    outputs(9729) <= layer2_outputs(2668);
    outputs(9730) <= not(layer2_outputs(8019));
    outputs(9731) <= not(layer2_outputs(5321)) or (layer2_outputs(5866));
    outputs(9732) <= not(layer2_outputs(497));
    outputs(9733) <= layer2_outputs(53);
    outputs(9734) <= layer2_outputs(2909);
    outputs(9735) <= not(layer2_outputs(1054));
    outputs(9736) <= (layer2_outputs(457)) and not (layer2_outputs(8962));
    outputs(9737) <= not((layer2_outputs(6358)) xor (layer2_outputs(135)));
    outputs(9738) <= not(layer2_outputs(6707));
    outputs(9739) <= (layer2_outputs(4051)) and not (layer2_outputs(1072));
    outputs(9740) <= not(layer2_outputs(8219));
    outputs(9741) <= layer2_outputs(6990);
    outputs(9742) <= not(layer2_outputs(8063)) or (layer2_outputs(8071));
    outputs(9743) <= not((layer2_outputs(1661)) xor (layer2_outputs(3357)));
    outputs(9744) <= layer2_outputs(4945);
    outputs(9745) <= (layer2_outputs(8892)) and not (layer2_outputs(6516));
    outputs(9746) <= not(layer2_outputs(6619));
    outputs(9747) <= (layer2_outputs(1082)) and not (layer2_outputs(5168));
    outputs(9748) <= not(layer2_outputs(4885)) or (layer2_outputs(8662));
    outputs(9749) <= layer2_outputs(8444);
    outputs(9750) <= layer2_outputs(1723);
    outputs(9751) <= layer2_outputs(6856);
    outputs(9752) <= not((layer2_outputs(3470)) or (layer2_outputs(6952)));
    outputs(9753) <= not(layer2_outputs(9339));
    outputs(9754) <= not((layer2_outputs(6499)) xor (layer2_outputs(6246)));
    outputs(9755) <= layer2_outputs(538);
    outputs(9756) <= (layer2_outputs(3249)) and not (layer2_outputs(2009));
    outputs(9757) <= not((layer2_outputs(9111)) or (layer2_outputs(345)));
    outputs(9758) <= layer2_outputs(1849);
    outputs(9759) <= not((layer2_outputs(7821)) and (layer2_outputs(7225)));
    outputs(9760) <= not(layer2_outputs(1323));
    outputs(9761) <= not((layer2_outputs(412)) and (layer2_outputs(3354)));
    outputs(9762) <= not(layer2_outputs(3766)) or (layer2_outputs(8069));
    outputs(9763) <= not(layer2_outputs(762)) or (layer2_outputs(6827));
    outputs(9764) <= not((layer2_outputs(5756)) xor (layer2_outputs(5628)));
    outputs(9765) <= not(layer2_outputs(4163));
    outputs(9766) <= not(layer2_outputs(10052));
    outputs(9767) <= not(layer2_outputs(4646));
    outputs(9768) <= not(layer2_outputs(2855));
    outputs(9769) <= not((layer2_outputs(683)) xor (layer2_outputs(4874)));
    outputs(9770) <= (layer2_outputs(1984)) xor (layer2_outputs(4455));
    outputs(9771) <= (layer2_outputs(4275)) and not (layer2_outputs(3241));
    outputs(9772) <= (layer2_outputs(480)) and not (layer2_outputs(6206));
    outputs(9773) <= not(layer2_outputs(7509));
    outputs(9774) <= not(layer2_outputs(2856));
    outputs(9775) <= (layer2_outputs(4101)) xor (layer2_outputs(6137));
    outputs(9776) <= not(layer2_outputs(9360));
    outputs(9777) <= not(layer2_outputs(9610));
    outputs(9778) <= not(layer2_outputs(7801));
    outputs(9779) <= layer2_outputs(3558);
    outputs(9780) <= layer2_outputs(3258);
    outputs(9781) <= layer2_outputs(5229);
    outputs(9782) <= layer2_outputs(2967);
    outputs(9783) <= not(layer2_outputs(7749));
    outputs(9784) <= not(layer2_outputs(7164));
    outputs(9785) <= not(layer2_outputs(7975));
    outputs(9786) <= (layer2_outputs(1056)) and (layer2_outputs(7269));
    outputs(9787) <= not(layer2_outputs(4565));
    outputs(9788) <= layer2_outputs(7000);
    outputs(9789) <= not(layer2_outputs(10035)) or (layer2_outputs(7026));
    outputs(9790) <= not((layer2_outputs(4442)) or (layer2_outputs(1324)));
    outputs(9791) <= not((layer2_outputs(1817)) xor (layer2_outputs(8932)));
    outputs(9792) <= not((layer2_outputs(2005)) and (layer2_outputs(5964)));
    outputs(9793) <= not(layer2_outputs(6703));
    outputs(9794) <= layer2_outputs(5672);
    outputs(9795) <= (layer2_outputs(1490)) and not (layer2_outputs(724));
    outputs(9796) <= not(layer2_outputs(4774));
    outputs(9797) <= not(layer2_outputs(1086)) or (layer2_outputs(2341));
    outputs(9798) <= not(layer2_outputs(9316));
    outputs(9799) <= (layer2_outputs(945)) xor (layer2_outputs(900));
    outputs(9800) <= not(layer2_outputs(8976));
    outputs(9801) <= layer2_outputs(105);
    outputs(9802) <= not(layer2_outputs(1950));
    outputs(9803) <= not(layer2_outputs(2064));
    outputs(9804) <= layer2_outputs(1061);
    outputs(9805) <= not(layer2_outputs(2904));
    outputs(9806) <= layer2_outputs(4472);
    outputs(9807) <= layer2_outputs(3206);
    outputs(9808) <= layer2_outputs(4331);
    outputs(9809) <= not(layer2_outputs(9840));
    outputs(9810) <= layer2_outputs(5895);
    outputs(9811) <= not(layer2_outputs(9830));
    outputs(9812) <= not(layer2_outputs(1154)) or (layer2_outputs(4512));
    outputs(9813) <= not(layer2_outputs(9970));
    outputs(9814) <= not(layer2_outputs(2325));
    outputs(9815) <= not((layer2_outputs(9819)) xor (layer2_outputs(931)));
    outputs(9816) <= not(layer2_outputs(9583));
    outputs(9817) <= not(layer2_outputs(4267));
    outputs(9818) <= layer2_outputs(5015);
    outputs(9819) <= not(layer2_outputs(1370));
    outputs(9820) <= not(layer2_outputs(8720));
    outputs(9821) <= not(layer2_outputs(2486));
    outputs(9822) <= not(layer2_outputs(650));
    outputs(9823) <= not((layer2_outputs(97)) xor (layer2_outputs(4894)));
    outputs(9824) <= layer2_outputs(3711);
    outputs(9825) <= not(layer2_outputs(8527));
    outputs(9826) <= not(layer2_outputs(2352));
    outputs(9827) <= layer2_outputs(3833);
    outputs(9828) <= not((layer2_outputs(10237)) or (layer2_outputs(9142)));
    outputs(9829) <= not((layer2_outputs(1494)) xor (layer2_outputs(4950)));
    outputs(9830) <= not((layer2_outputs(6342)) xor (layer2_outputs(5017)));
    outputs(9831) <= (layer2_outputs(4138)) xor (layer2_outputs(3376));
    outputs(9832) <= (layer2_outputs(8761)) xor (layer2_outputs(6940));
    outputs(9833) <= not((layer2_outputs(4224)) xor (layer2_outputs(5241)));
    outputs(9834) <= (layer2_outputs(20)) or (layer2_outputs(5245));
    outputs(9835) <= (layer2_outputs(2523)) and not (layer2_outputs(5699));
    outputs(9836) <= (layer2_outputs(2291)) xor (layer2_outputs(3281));
    outputs(9837) <= (layer2_outputs(2995)) and not (layer2_outputs(1848));
    outputs(9838) <= not((layer2_outputs(3734)) and (layer2_outputs(6312)));
    outputs(9839) <= (layer2_outputs(1763)) xor (layer2_outputs(335));
    outputs(9840) <= not(layer2_outputs(5486));
    outputs(9841) <= (layer2_outputs(3114)) and (layer2_outputs(5573));
    outputs(9842) <= not(layer2_outputs(6391));
    outputs(9843) <= (layer2_outputs(6793)) and not (layer2_outputs(880));
    outputs(9844) <= not(layer2_outputs(1204));
    outputs(9845) <= (layer2_outputs(186)) or (layer2_outputs(2358));
    outputs(9846) <= not((layer2_outputs(8568)) xor (layer2_outputs(1188)));
    outputs(9847) <= layer2_outputs(2834);
    outputs(9848) <= (layer2_outputs(3195)) xor (layer2_outputs(3356));
    outputs(9849) <= not(layer2_outputs(2966));
    outputs(9850) <= layer2_outputs(6679);
    outputs(9851) <= not((layer2_outputs(5705)) and (layer2_outputs(3306)));
    outputs(9852) <= layer2_outputs(86);
    outputs(9853) <= not((layer2_outputs(5759)) xor (layer2_outputs(5725)));
    outputs(9854) <= layer2_outputs(5735);
    outputs(9855) <= (layer2_outputs(5426)) and not (layer2_outputs(5341));
    outputs(9856) <= layer2_outputs(2847);
    outputs(9857) <= (layer2_outputs(2992)) and not (layer2_outputs(9815));
    outputs(9858) <= (layer2_outputs(6618)) and not (layer2_outputs(7499));
    outputs(9859) <= not(layer2_outputs(7371));
    outputs(9860) <= not(layer2_outputs(7284));
    outputs(9861) <= layer2_outputs(3521);
    outputs(9862) <= (layer2_outputs(8994)) and not (layer2_outputs(773));
    outputs(9863) <= not((layer2_outputs(4493)) xor (layer2_outputs(9858)));
    outputs(9864) <= not((layer2_outputs(5128)) xor (layer2_outputs(4348)));
    outputs(9865) <= not(layer2_outputs(6991));
    outputs(9866) <= layer2_outputs(4269);
    outputs(9867) <= layer2_outputs(7040);
    outputs(9868) <= not(layer2_outputs(373));
    outputs(9869) <= (layer2_outputs(7957)) and not (layer2_outputs(4392));
    outputs(9870) <= (layer2_outputs(2661)) and (layer2_outputs(6368));
    outputs(9871) <= not(layer2_outputs(3907));
    outputs(9872) <= layer2_outputs(845);
    outputs(9873) <= not(layer2_outputs(8379));
    outputs(9874) <= layer2_outputs(5707);
    outputs(9875) <= not((layer2_outputs(8686)) and (layer2_outputs(3807)));
    outputs(9876) <= not(layer2_outputs(461)) or (layer2_outputs(1909));
    outputs(9877) <= layer2_outputs(8170);
    outputs(9878) <= layer2_outputs(3680);
    outputs(9879) <= (layer2_outputs(5616)) xor (layer2_outputs(4423));
    outputs(9880) <= not(layer2_outputs(4600));
    outputs(9881) <= (layer2_outputs(5512)) and (layer2_outputs(4713));
    outputs(9882) <= layer2_outputs(3990);
    outputs(9883) <= not(layer2_outputs(1945));
    outputs(9884) <= layer2_outputs(1065);
    outputs(9885) <= (layer2_outputs(6930)) xor (layer2_outputs(1782));
    outputs(9886) <= (layer2_outputs(2051)) and not (layer2_outputs(8847));
    outputs(9887) <= layer2_outputs(7622);
    outputs(9888) <= (layer2_outputs(4177)) xor (layer2_outputs(8264));
    outputs(9889) <= layer2_outputs(7716);
    outputs(9890) <= not((layer2_outputs(2622)) xor (layer2_outputs(6423)));
    outputs(9891) <= (layer2_outputs(3225)) and (layer2_outputs(5166));
    outputs(9892) <= (layer2_outputs(5246)) and not (layer2_outputs(6544));
    outputs(9893) <= layer2_outputs(612);
    outputs(9894) <= (layer2_outputs(350)) xor (layer2_outputs(7633));
    outputs(9895) <= not(layer2_outputs(2916));
    outputs(9896) <= not(layer2_outputs(9997));
    outputs(9897) <= layer2_outputs(8667);
    outputs(9898) <= layer2_outputs(8547);
    outputs(9899) <= not(layer2_outputs(1961)) or (layer2_outputs(5318));
    outputs(9900) <= not(layer2_outputs(4082)) or (layer2_outputs(7365));
    outputs(9901) <= (layer2_outputs(2565)) xor (layer2_outputs(8422));
    outputs(9902) <= layer2_outputs(4420);
    outputs(9903) <= not(layer2_outputs(7637));
    outputs(9904) <= layer2_outputs(8526);
    outputs(9905) <= not((layer2_outputs(4362)) xor (layer2_outputs(57)));
    outputs(9906) <= (layer2_outputs(2678)) xor (layer2_outputs(3685));
    outputs(9907) <= not(layer2_outputs(3658));
    outputs(9908) <= not((layer2_outputs(1540)) or (layer2_outputs(1700)));
    outputs(9909) <= (layer2_outputs(2948)) xor (layer2_outputs(6035));
    outputs(9910) <= not(layer2_outputs(720));
    outputs(9911) <= (layer2_outputs(2369)) and (layer2_outputs(3207));
    outputs(9912) <= layer2_outputs(8038);
    outputs(9913) <= layer2_outputs(2461);
    outputs(9914) <= not(layer2_outputs(4118));
    outputs(9915) <= not(layer2_outputs(1717));
    outputs(9916) <= not((layer2_outputs(5072)) xor (layer2_outputs(9088)));
    outputs(9917) <= not((layer2_outputs(3168)) xor (layer2_outputs(469)));
    outputs(9918) <= layer2_outputs(4088);
    outputs(9919) <= (layer2_outputs(2901)) xor (layer2_outputs(5359));
    outputs(9920) <= not(layer2_outputs(5696));
    outputs(9921) <= layer2_outputs(6060);
    outputs(9922) <= layer2_outputs(3545);
    outputs(9923) <= (layer2_outputs(3526)) or (layer2_outputs(9994));
    outputs(9924) <= layer2_outputs(7512);
    outputs(9925) <= not((layer2_outputs(1529)) xor (layer2_outputs(6725)));
    outputs(9926) <= (layer2_outputs(5347)) xor (layer2_outputs(2217));
    outputs(9927) <= (layer2_outputs(7680)) and (layer2_outputs(2330));
    outputs(9928) <= layer2_outputs(976);
    outputs(9929) <= layer2_outputs(5739);
    outputs(9930) <= not((layer2_outputs(7213)) and (layer2_outputs(10200)));
    outputs(9931) <= not(layer2_outputs(9333)) or (layer2_outputs(8392));
    outputs(9932) <= not((layer2_outputs(10091)) or (layer2_outputs(935)));
    outputs(9933) <= (layer2_outputs(6011)) and not (layer2_outputs(3629));
    outputs(9934) <= not(layer2_outputs(3962));
    outputs(9935) <= not(layer2_outputs(2552));
    outputs(9936) <= layer2_outputs(8369);
    outputs(9937) <= not(layer2_outputs(2582));
    outputs(9938) <= layer2_outputs(1001);
    outputs(9939) <= not(layer2_outputs(9630));
    outputs(9940) <= (layer2_outputs(7919)) and not (layer2_outputs(4087));
    outputs(9941) <= not((layer2_outputs(3307)) xor (layer2_outputs(3569)));
    outputs(9942) <= (layer2_outputs(7482)) xor (layer2_outputs(8788));
    outputs(9943) <= (layer2_outputs(5402)) xor (layer2_outputs(7161));
    outputs(9944) <= layer2_outputs(4012);
    outputs(9945) <= not((layer2_outputs(8436)) xor (layer2_outputs(753)));
    outputs(9946) <= (layer2_outputs(3941)) and (layer2_outputs(9138));
    outputs(9947) <= (layer2_outputs(270)) and not (layer2_outputs(7760));
    outputs(9948) <= layer2_outputs(9939);
    outputs(9949) <= not(layer2_outputs(2437));
    outputs(9950) <= (layer2_outputs(2077)) xor (layer2_outputs(2881));
    outputs(9951) <= layer2_outputs(10115);
    outputs(9952) <= (layer2_outputs(6645)) xor (layer2_outputs(3029));
    outputs(9953) <= not((layer2_outputs(5287)) xor (layer2_outputs(9174)));
    outputs(9954) <= not(layer2_outputs(681));
    outputs(9955) <= not(layer2_outputs(6789));
    outputs(9956) <= (layer2_outputs(8100)) xor (layer2_outputs(7855));
    outputs(9957) <= layer2_outputs(3233);
    outputs(9958) <= not((layer2_outputs(5860)) xor (layer2_outputs(5273)));
    outputs(9959) <= not(layer2_outputs(964));
    outputs(9960) <= layer2_outputs(2562);
    outputs(9961) <= (layer2_outputs(324)) or (layer2_outputs(9260));
    outputs(9962) <= (layer2_outputs(5822)) and not (layer2_outputs(3142));
    outputs(9963) <= layer2_outputs(1608);
    outputs(9964) <= not(layer2_outputs(6053));
    outputs(9965) <= (layer2_outputs(893)) and not (layer2_outputs(4758));
    outputs(9966) <= not(layer2_outputs(8057));
    outputs(9967) <= not(layer2_outputs(2848));
    outputs(9968) <= not(layer2_outputs(10071));
    outputs(9969) <= not((layer2_outputs(1214)) xor (layer2_outputs(191)));
    outputs(9970) <= not((layer2_outputs(10073)) or (layer2_outputs(6643)));
    outputs(9971) <= not(layer2_outputs(3741));
    outputs(9972) <= layer2_outputs(274);
    outputs(9973) <= layer2_outputs(5155);
    outputs(9974) <= layer2_outputs(271);
    outputs(9975) <= not(layer2_outputs(7182)) or (layer2_outputs(9694));
    outputs(9976) <= not(layer2_outputs(2966));
    outputs(9977) <= layer2_outputs(9493);
    outputs(9978) <= (layer2_outputs(837)) and not (layer2_outputs(3535));
    outputs(9979) <= not(layer2_outputs(187));
    outputs(9980) <= not(layer2_outputs(5055));
    outputs(9981) <= not(layer2_outputs(4267));
    outputs(9982) <= not(layer2_outputs(2057));
    outputs(9983) <= not(layer2_outputs(6519)) or (layer2_outputs(3283));
    outputs(9984) <= layer2_outputs(1886);
    outputs(9985) <= layer2_outputs(6493);
    outputs(9986) <= not((layer2_outputs(9202)) or (layer2_outputs(90)));
    outputs(9987) <= not(layer2_outputs(475));
    outputs(9988) <= not((layer2_outputs(9833)) xor (layer2_outputs(9600)));
    outputs(9989) <= not(layer2_outputs(3695));
    outputs(9990) <= not(layer2_outputs(7857)) or (layer2_outputs(10016));
    outputs(9991) <= not((layer2_outputs(622)) or (layer2_outputs(5681)));
    outputs(9992) <= not(layer2_outputs(772));
    outputs(9993) <= not((layer2_outputs(2273)) and (layer2_outputs(9393)));
    outputs(9994) <= (layer2_outputs(10094)) xor (layer2_outputs(8184));
    outputs(9995) <= not((layer2_outputs(7403)) xor (layer2_outputs(8081)));
    outputs(9996) <= (layer2_outputs(3897)) and not (layer2_outputs(8829));
    outputs(9997) <= not(layer2_outputs(9564));
    outputs(9998) <= not(layer2_outputs(5308));
    outputs(9999) <= (layer2_outputs(2718)) and (layer2_outputs(9295));
    outputs(10000) <= not(layer2_outputs(9554));
    outputs(10001) <= not(layer2_outputs(956)) or (layer2_outputs(8052));
    outputs(10002) <= not(layer2_outputs(2741));
    outputs(10003) <= (layer2_outputs(4073)) and (layer2_outputs(7324));
    outputs(10004) <= not((layer2_outputs(10198)) xor (layer2_outputs(9097)));
    outputs(10005) <= (layer2_outputs(3422)) and (layer2_outputs(3738));
    outputs(10006) <= layer2_outputs(4837);
    outputs(10007) <= (layer2_outputs(1372)) xor (layer2_outputs(6840));
    outputs(10008) <= not(layer2_outputs(4105));
    outputs(10009) <= not(layer2_outputs(1111));
    outputs(10010) <= (layer2_outputs(7562)) xor (layer2_outputs(4013));
    outputs(10011) <= not(layer2_outputs(6868)) or (layer2_outputs(9222));
    outputs(10012) <= (layer2_outputs(537)) xor (layer2_outputs(676));
    outputs(10013) <= layer2_outputs(1432);
    outputs(10014) <= not(layer2_outputs(8665));
    outputs(10015) <= not(layer2_outputs(4842));
    outputs(10016) <= not((layer2_outputs(7470)) xor (layer2_outputs(4814)));
    outputs(10017) <= layer2_outputs(4756);
    outputs(10018) <= layer2_outputs(3025);
    outputs(10019) <= layer2_outputs(8210);
    outputs(10020) <= not((layer2_outputs(529)) xor (layer2_outputs(8842)));
    outputs(10021) <= layer2_outputs(9924);
    outputs(10022) <= (layer2_outputs(3714)) or (layer2_outputs(3088));
    outputs(10023) <= not(layer2_outputs(8229));
    outputs(10024) <= layer2_outputs(1056);
    outputs(10025) <= layer2_outputs(6967);
    outputs(10026) <= layer2_outputs(7805);
    outputs(10027) <= (layer2_outputs(3463)) xor (layer2_outputs(2685));
    outputs(10028) <= not(layer2_outputs(5593));
    outputs(10029) <= layer2_outputs(6823);
    outputs(10030) <= (layer2_outputs(4935)) and not (layer2_outputs(2555));
    outputs(10031) <= not(layer2_outputs(2907));
    outputs(10032) <= not((layer2_outputs(531)) xor (layer2_outputs(3628)));
    outputs(10033) <= not((layer2_outputs(6346)) xor (layer2_outputs(9807)));
    outputs(10034) <= layer2_outputs(2386);
    outputs(10035) <= layer2_outputs(8662);
    outputs(10036) <= layer2_outputs(7234);
    outputs(10037) <= not(layer2_outputs(6020));
    outputs(10038) <= '0';
    outputs(10039) <= layer2_outputs(2417);
    outputs(10040) <= not((layer2_outputs(8415)) and (layer2_outputs(7408)));
    outputs(10041) <= layer2_outputs(348);
    outputs(10042) <= not((layer2_outputs(3153)) xor (layer2_outputs(7059)));
    outputs(10043) <= not(layer2_outputs(8792)) or (layer2_outputs(5416));
    outputs(10044) <= (layer2_outputs(5893)) xor (layer2_outputs(5871));
    outputs(10045) <= not(layer2_outputs(5097)) or (layer2_outputs(580));
    outputs(10046) <= not((layer2_outputs(6130)) or (layer2_outputs(5700)));
    outputs(10047) <= not(layer2_outputs(9066));
    outputs(10048) <= layer2_outputs(9835);
    outputs(10049) <= (layer2_outputs(5885)) and not (layer2_outputs(2036));
    outputs(10050) <= (layer2_outputs(4047)) xor (layer2_outputs(5252));
    outputs(10051) <= not(layer2_outputs(635));
    outputs(10052) <= not(layer2_outputs(9923));
    outputs(10053) <= not(layer2_outputs(229));
    outputs(10054) <= layer2_outputs(3820);
    outputs(10055) <= (layer2_outputs(6673)) or (layer2_outputs(8978));
    outputs(10056) <= layer2_outputs(6110);
    outputs(10057) <= not((layer2_outputs(1044)) or (layer2_outputs(3397)));
    outputs(10058) <= layer2_outputs(10238);
    outputs(10059) <= (layer2_outputs(7668)) xor (layer2_outputs(164));
    outputs(10060) <= not((layer2_outputs(7840)) xor (layer2_outputs(1776)));
    outputs(10061) <= (layer2_outputs(2896)) xor (layer2_outputs(209));
    outputs(10062) <= not(layer2_outputs(7394));
    outputs(10063) <= not((layer2_outputs(4394)) xor (layer2_outputs(6111)));
    outputs(10064) <= layer2_outputs(6804);
    outputs(10065) <= not(layer2_outputs(8036));
    outputs(10066) <= (layer2_outputs(9176)) xor (layer2_outputs(3311));
    outputs(10067) <= (layer2_outputs(4279)) xor (layer2_outputs(1233));
    outputs(10068) <= layer2_outputs(9107);
    outputs(10069) <= layer2_outputs(4738);
    outputs(10070) <= layer2_outputs(9953);
    outputs(10071) <= not(layer2_outputs(8504));
    outputs(10072) <= not((layer2_outputs(750)) xor (layer2_outputs(2538)));
    outputs(10073) <= (layer2_outputs(3391)) and not (layer2_outputs(8223));
    outputs(10074) <= (layer2_outputs(8622)) and (layer2_outputs(2408));
    outputs(10075) <= layer2_outputs(2509);
    outputs(10076) <= not(layer2_outputs(8602));
    outputs(10077) <= not((layer2_outputs(2413)) and (layer2_outputs(8423)));
    outputs(10078) <= layer2_outputs(2114);
    outputs(10079) <= layer2_outputs(4397);
    outputs(10080) <= not(layer2_outputs(3693)) or (layer2_outputs(5181));
    outputs(10081) <= not((layer2_outputs(9119)) xor (layer2_outputs(4846)));
    outputs(10082) <= layer2_outputs(1726);
    outputs(10083) <= not((layer2_outputs(9031)) xor (layer2_outputs(5202)));
    outputs(10084) <= layer2_outputs(3094);
    outputs(10085) <= (layer2_outputs(5159)) and not (layer2_outputs(4217));
    outputs(10086) <= (layer2_outputs(8999)) xor (layer2_outputs(8328));
    outputs(10087) <= (layer2_outputs(5927)) xor (layer2_outputs(7836));
    outputs(10088) <= layer2_outputs(1205);
    outputs(10089) <= layer2_outputs(2758);
    outputs(10090) <= not((layer2_outputs(7802)) xor (layer2_outputs(498)));
    outputs(10091) <= layer2_outputs(9526);
    outputs(10092) <= (layer2_outputs(9908)) xor (layer2_outputs(7391));
    outputs(10093) <= layer2_outputs(1428);
    outputs(10094) <= not((layer2_outputs(1052)) xor (layer2_outputs(8718)));
    outputs(10095) <= layer2_outputs(6906);
    outputs(10096) <= layer2_outputs(3245);
    outputs(10097) <= not((layer2_outputs(437)) xor (layer2_outputs(7600)));
    outputs(10098) <= not(layer2_outputs(4995));
    outputs(10099) <= not(layer2_outputs(8513));
    outputs(10100) <= (layer2_outputs(5084)) xor (layer2_outputs(9366));
    outputs(10101) <= (layer2_outputs(8475)) xor (layer2_outputs(9649));
    outputs(10102) <= (layer2_outputs(2054)) xor (layer2_outputs(7900));
    outputs(10103) <= (layer2_outputs(4994)) and not (layer2_outputs(1766));
    outputs(10104) <= not((layer2_outputs(8888)) or (layer2_outputs(5023)));
    outputs(10105) <= not((layer2_outputs(543)) xor (layer2_outputs(7494)));
    outputs(10106) <= (layer2_outputs(3499)) and (layer2_outputs(4301));
    outputs(10107) <= not(layer2_outputs(3438));
    outputs(10108) <= (layer2_outputs(1018)) or (layer2_outputs(5840));
    outputs(10109) <= layer2_outputs(655);
    outputs(10110) <= (layer2_outputs(7559)) and not (layer2_outputs(4750));
    outputs(10111) <= (layer2_outputs(979)) xor (layer2_outputs(5809));
    outputs(10112) <= (layer2_outputs(1028)) xor (layer2_outputs(3265));
    outputs(10113) <= not(layer2_outputs(7337));
    outputs(10114) <= not(layer2_outputs(9726));
    outputs(10115) <= not(layer2_outputs(500));
    outputs(10116) <= not((layer2_outputs(633)) xor (layer2_outputs(8730)));
    outputs(10117) <= not(layer2_outputs(9273));
    outputs(10118) <= (layer2_outputs(9688)) or (layer2_outputs(6508));
    outputs(10119) <= layer2_outputs(53);
    outputs(10120) <= (layer2_outputs(8256)) and not (layer2_outputs(6146));
    outputs(10121) <= not((layer2_outputs(7394)) or (layer2_outputs(1583)));
    outputs(10122) <= layer2_outputs(10097);
    outputs(10123) <= not(layer2_outputs(2743));
    outputs(10124) <= not((layer2_outputs(10215)) or (layer2_outputs(5119)));
    outputs(10125) <= not((layer2_outputs(6123)) xor (layer2_outputs(932)));
    outputs(10126) <= layer2_outputs(7678);
    outputs(10127) <= not(layer2_outputs(8357));
    outputs(10128) <= not(layer2_outputs(1545));
    outputs(10129) <= not((layer2_outputs(9878)) xor (layer2_outputs(9798)));
    outputs(10130) <= (layer2_outputs(3627)) and not (layer2_outputs(8074));
    outputs(10131) <= (layer2_outputs(7243)) or (layer2_outputs(6834));
    outputs(10132) <= not(layer2_outputs(2241));
    outputs(10133) <= layer2_outputs(3729);
    outputs(10134) <= not((layer2_outputs(4166)) xor (layer2_outputs(5169)));
    outputs(10135) <= layer2_outputs(8530);
    outputs(10136) <= not(layer2_outputs(6176)) or (layer2_outputs(9281));
    outputs(10137) <= not((layer2_outputs(4313)) or (layer2_outputs(9326)));
    outputs(10138) <= not(layer2_outputs(7424));
    outputs(10139) <= '1';
    outputs(10140) <= not(layer2_outputs(9358));
    outputs(10141) <= layer2_outputs(5910);
    outputs(10142) <= not((layer2_outputs(1529)) or (layer2_outputs(4329)));
    outputs(10143) <= layer2_outputs(5404);
    outputs(10144) <= layer2_outputs(465);
    outputs(10145) <= not((layer2_outputs(2138)) xor (layer2_outputs(4494)));
    outputs(10146) <= not((layer2_outputs(157)) xor (layer2_outputs(8777)));
    outputs(10147) <= not(layer2_outputs(4146));
    outputs(10148) <= (layer2_outputs(7909)) and not (layer2_outputs(467));
    outputs(10149) <= layer2_outputs(5014);
    outputs(10150) <= not(layer2_outputs(343));
    outputs(10151) <= not(layer2_outputs(9873));
    outputs(10152) <= layer2_outputs(9246);
    outputs(10153) <= not(layer2_outputs(8516));
    outputs(10154) <= (layer2_outputs(4245)) xor (layer2_outputs(8307));
    outputs(10155) <= not(layer2_outputs(4294));
    outputs(10156) <= layer2_outputs(7413);
    outputs(10157) <= layer2_outputs(543);
    outputs(10158) <= not((layer2_outputs(3064)) xor (layer2_outputs(8938)));
    outputs(10159) <= layer2_outputs(5146);
    outputs(10160) <= not((layer2_outputs(7017)) xor (layer2_outputs(9468)));
    outputs(10161) <= not(layer2_outputs(6156));
    outputs(10162) <= not((layer2_outputs(7971)) xor (layer2_outputs(1407)));
    outputs(10163) <= not(layer2_outputs(9287));
    outputs(10164) <= (layer2_outputs(8776)) and not (layer2_outputs(2835));
    outputs(10165) <= (layer2_outputs(8425)) and not (layer2_outputs(7938));
    outputs(10166) <= not(layer2_outputs(8717));
    outputs(10167) <= not(layer2_outputs(10205));
    outputs(10168) <= not(layer2_outputs(2841));
    outputs(10169) <= not(layer2_outputs(7536));
    outputs(10170) <= not(layer2_outputs(7947));
    outputs(10171) <= not(layer2_outputs(9811));
    outputs(10172) <= not(layer2_outputs(102));
    outputs(10173) <= (layer2_outputs(3601)) and (layer2_outputs(6593));
    outputs(10174) <= not(layer2_outputs(6763));
    outputs(10175) <= (layer2_outputs(4514)) and not (layer2_outputs(1401));
    outputs(10176) <= not(layer2_outputs(3178));
    outputs(10177) <= '1';
    outputs(10178) <= layer2_outputs(8523);
    outputs(10179) <= layer2_outputs(2299);
    outputs(10180) <= not(layer2_outputs(5524));
    outputs(10181) <= (layer2_outputs(4978)) and not (layer2_outputs(1261));
    outputs(10182) <= (layer2_outputs(1734)) xor (layer2_outputs(683));
    outputs(10183) <= not((layer2_outputs(3592)) xor (layer2_outputs(8959)));
    outputs(10184) <= (layer2_outputs(6038)) xor (layer2_outputs(8272));
    outputs(10185) <= layer2_outputs(4460);
    outputs(10186) <= not(layer2_outputs(7646));
    outputs(10187) <= layer2_outputs(8260);
    outputs(10188) <= (layer2_outputs(9991)) and not (layer2_outputs(9082));
    outputs(10189) <= not(layer2_outputs(3057));
    outputs(10190) <= (layer2_outputs(9561)) and not (layer2_outputs(4989));
    outputs(10191) <= (layer2_outputs(4726)) and (layer2_outputs(4790));
    outputs(10192) <= layer2_outputs(1842);
    outputs(10193) <= layer2_outputs(1033);
    outputs(10194) <= (layer2_outputs(7892)) and not (layer2_outputs(8772));
    outputs(10195) <= (layer2_outputs(344)) xor (layer2_outputs(7377));
    outputs(10196) <= layer2_outputs(1451);
    outputs(10197) <= (layer2_outputs(1493)) xor (layer2_outputs(2152));
    outputs(10198) <= layer2_outputs(7429);
    outputs(10199) <= (layer2_outputs(5967)) xor (layer2_outputs(646));
    outputs(10200) <= not((layer2_outputs(4626)) and (layer2_outputs(3093)));
    outputs(10201) <= not(layer2_outputs(1879));
    outputs(10202) <= layer2_outputs(2987);
    outputs(10203) <= not(layer2_outputs(7505));
    outputs(10204) <= not(layer2_outputs(1484));
    outputs(10205) <= not((layer2_outputs(6042)) and (layer2_outputs(1372)));
    outputs(10206) <= layer2_outputs(8889);
    outputs(10207) <= not((layer2_outputs(8991)) or (layer2_outputs(2087)));
    outputs(10208) <= layer2_outputs(9321);
    outputs(10209) <= not(layer2_outputs(6999));
    outputs(10210) <= not(layer2_outputs(2263));
    outputs(10211) <= layer2_outputs(7931);
    outputs(10212) <= not(layer2_outputs(758));
    outputs(10213) <= not(layer2_outputs(8686));
    outputs(10214) <= not(layer2_outputs(1963));
    outputs(10215) <= (layer2_outputs(9394)) and not (layer2_outputs(1449));
    outputs(10216) <= (layer2_outputs(5130)) and (layer2_outputs(3276));
    outputs(10217) <= (layer2_outputs(1413)) and (layer2_outputs(5605));
    outputs(10218) <= (layer2_outputs(9345)) and not (layer2_outputs(7874));
    outputs(10219) <= layer2_outputs(10101);
    outputs(10220) <= not(layer2_outputs(8838));
    outputs(10221) <= (layer2_outputs(6074)) or (layer2_outputs(3146));
    outputs(10222) <= not(layer2_outputs(9883));
    outputs(10223) <= layer2_outputs(3514);
    outputs(10224) <= not((layer2_outputs(4916)) xor (layer2_outputs(5677)));
    outputs(10225) <= (layer2_outputs(49)) xor (layer2_outputs(358));
    outputs(10226) <= (layer2_outputs(2299)) and not (layer2_outputs(5297));
    outputs(10227) <= layer2_outputs(5335);
    outputs(10228) <= (layer2_outputs(1615)) xor (layer2_outputs(571));
    outputs(10229) <= layer2_outputs(6634);
    outputs(10230) <= layer2_outputs(51);
    outputs(10231) <= not(layer2_outputs(3718));
    outputs(10232) <= not(layer2_outputs(7950));
    outputs(10233) <= not(layer2_outputs(4850));
    outputs(10234) <= (layer2_outputs(952)) xor (layer2_outputs(2067));
    outputs(10235) <= not(layer2_outputs(1300));
    outputs(10236) <= layer2_outputs(1230);
    outputs(10237) <= not((layer2_outputs(6505)) and (layer2_outputs(10009)));
    outputs(10238) <= layer2_outputs(6526);
    outputs(10239) <= layer2_outputs(2110);

end Behavioral;
